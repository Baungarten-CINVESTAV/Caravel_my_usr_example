* NGSPICE file created from m_Top_Module_User.ext - technology: sky130B

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR Y B1 A2 A1 A3 VNB VPB
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_1 C B Y D A VPWR VGND VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41oi_4 B1 A2 A1 A4 A3 Y VGND VPWR VNB VPB
X0 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A1 a_493_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A4 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A1 a_493_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_911_47# A2 a_493_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_911_47# A3 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A4 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A4 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_493_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_493_47# A2 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_493_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_493_47# A2 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_911_47# A2 a_493_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_1269_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_911_47# A3 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_27_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VPWR A4 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_1269_47# A3 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_27_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_1269_47# A3 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_1269_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR B X A_N C VNB VPB
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_4 B C A D X VPWR VGND VNB VPB
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A X VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_1 A2 B1 A1 A3 X VGND VPWR VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N X A2_N B2 B1 VPWR VGND VNB VPB
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_1 Y A C B VGND VPWR VNB VPB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND A X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_4 Y B1 A2 A1 VPWR VGND VNB VPB
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4b_2 D C B Y A_N VGND VPWR VNB VPB
X0 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_465_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND D a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_215_47# B a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_655_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_655_47# C a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_465_47# C a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR VNB VPB
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_1 Y A1_N A2_N B2 B1 VGND VPWR VNB VPB
X0 VPWR A2_N a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y a_112_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B2 a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_297# A2_N a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_112_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_112_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR B1 a_478_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_394_47# a_112_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_394_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_478_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4b_4 D C B Y A_N VGND VPWR VNB VPB
X0 a_991_47# C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_991_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_991_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND D a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND D a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_633_47# C a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_633_47# C a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_991_47# C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 Y A B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_1 B C A_N Y VGND VPWR VNB VPB
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_4 A D C B Y VPWR VGND VNB VPB
X0 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 B1 A2 A1 Y VGND VPWR VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VNB VPB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_1 A X B C VPWR VGND VNB VPB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 Y VGND VPWR VNB VPB
X0 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 B1 Y A2 VPWR VGND VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_4 A2 B2 A1 B1 Y VGND VPWR VNB VPB
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_4 A C Y D B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VNB VPB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_1 B1 A1 B2 A2 Y VPWR VGND VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311oi_4 Y B1 A1 A3 C1 A2 VPWR VGND VNB VPB
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1139_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_1139_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_109_297# B1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_1139_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y C1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1139_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y C1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_4 A_N Y B C VGND VPWR VNB VPB
X0 VGND C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_633_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_633_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N Y VGND VPWR B2 B1 A2_N VNB VPB
X0 a_109_47# A2_N a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_397_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2_N a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_397_297# a_109_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_481_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B1 a_481_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_1 C A X B D VPWR VGND VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3b_4 A_N X C B VGND VPWR VNB VPB
X0 a_98_199# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_98_199# a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_257_47# B a_152_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_152_47# a_98_199# a_56_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR C a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_98_199# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_56_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND C a_257_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_2 B A Y D C VGND VPWR VNB VPB
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VNB VPB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_2 VPWR VGND X B A_N VNB VPB
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 D1 C1 A2 A1 B1 Y VGND VPWR VNB VPB
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_1 X A2 B1 A1 A3 VGND VPWR VNB VPB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_1 A2 A1 B1 X VPWR VGND VNB VPB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 Y C1 B1 VGND VPWR VNB VPB
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_1 Y A2 A1 A3 B1 VPWR VGND VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VPWR VGND VNB VPB
X0 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_762_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_80_21# A2 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A1 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_934_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_2 B2 Y A1_N A2_N B1 VGND VPWR VNB VPB
X0 a_113_297# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_113_47# A2_N a_113_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A2_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_730_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_471_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_471_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B2 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_113_297# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_113_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A1_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_113_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_113_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y a_113_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_730_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y a_113_297# a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_471_47# a_113_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR A1_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4bb_4 D_N B A C_N X VGND VPWR VNB VPB
X0 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_315_380# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A a_583_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_410# a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_583_297# B a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_397_297# a_205_93# a_315_380# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_499_297# a_27_410# a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_315_380# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A X VGND VPWR VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_16 Y A VGND VPWR VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A X VGND VPWR VNB VPB
X0 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=500000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=500000u
X3 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X7 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_4 B A_N Y VGND VPWR VNB VPB
X0 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_2 A Y B C VGND VPWR VNB VPB
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_2 A3 B1 Y A1 A2 VPWR VGND VNB VPB
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A2 B1 Y A1 B2 VGND VPWR VNB VPB
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR A1 A0 S X VNB VPB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 Y VPWR VGND VNB VPB
X0 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_298_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_664_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_298_47# B1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_497_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_497_47# B1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A2 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_27_47# C1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_497_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A1 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_664_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_2 C A X B D VPWR VGND VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N B1 B2 A2_N Y VGND VPWR VNB VPB
X0 a_1241_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_113_47# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_807_47# a_113_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B2 a_807_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_113_47# A2_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B2 a_807_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A2_N a_113_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y a_113_47# a_807_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_1241_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y B2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y a_113_47# a_807_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_807_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A1_N a_113_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_113_47# A2_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_807_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_807_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_1241_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR a_113_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_27_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_807_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_113_47# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y B2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y a_113_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VPWR a_113_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_113_47# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1241_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND A1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND B1 a_807_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 Y a_113_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND A1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND B1 a_807_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR B1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR A1_N a_113_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_113_47# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR A2_N a_113_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_807_47# a_113_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N X VPWR VGND VNB VPB
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR C A_N X D B VNB VPB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt m_Top_Module_User VGND VPWR io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] irq[0] irq[1] irq[2] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XFILLER_171_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0717__A0 _1486_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_46_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input92_A wbs_dat_i[28] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0708__A0 _1010_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_83_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1444__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__0986__C _1050_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_hold3_A hold3/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_123_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1270_ _1478_/A _1166_/Y _1270_/D _1281_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_95_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0985_ VPWR VGND _1050_/B _0985_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_118_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1468_ VGND VPWR _1468_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_921 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1374__287 la_data_out[65] _1374__287/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_26_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1439__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_186_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0770_ VGND VPWR _0770_/S _1301_/Q _1125_/B _0771_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_139_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_692 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1322_ _1322_/Q hold1/X _1322_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_96_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1614 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1253_ VGND VPWR _1247_/X _1246_/X _1248_/X _1253_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_56_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1106__B1 _1105_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_49_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1184_ VGND VPWR _1180_/X _1179_/X _1181_/X _1184_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_0_1703 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0880__A2 _1142_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_59_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0968_ _0970_/A _0986_/A _0979_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_140_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0899_ VGND VPWR _0899_/Y _0898_/X _0889_/Y _0849_/A _0891_/B VGND VPWR sky130_fd_sc_hd__a31oi_1
XFILLER_31_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput220 VPWR VGND wbs_dat_o[17] _0693_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput231 VPWR VGND wbs_dat_o[27] _0640_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_160_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput242 VPWR VGND wbs_dat_o[8] _0741_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_118_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1084__A _1132_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_27_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0856__C1 _0855_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_83_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_740 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_401 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input55_A la_oenb[52] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_117_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_154 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output211_A _1298_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1169__A _1203_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_187_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0822_ _0822_/C _0822_/B _0875_/A _0822_/D _0822_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_70_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0753_ VGND VPWR _0767_/S _1102_/A _1305_/Q _0754_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_171_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0801__A _1489_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_50_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0684_ VGND VPWR _0689_/S _1493_/A _1318_/Q _0685_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_192_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1305_ _1305_/Q _1228_/Y _1305_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_57_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1236_ VGND VPWR _1231_/X _1230_/X _1232_/X _1236_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_42_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1167_ VGND VPWR _1160_/X _1158_/X _1162_/X _1167_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_52_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1098_ _1097_/Y _1067_/A _1088_/X _1096_/Y _1093_/Y _1273_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41oi_4
XFILLER_52_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_743 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1079__A _1079_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1315__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0844__A2 input96/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_182_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_703 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output161_A _1496_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_136_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1452__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1430__343 la_data_out[121] _1430__343/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_94_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1021_ VGND VPWR _1021_/B _1021_/X _0813_/C _1021_/C VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_47_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0805_ _0805_/B _0838_/D _0805_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_50_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0736_ VGND VPWR _0742_/S _1059_/B _1308_/Q _0737_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_157_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0667_ VPWR VGND _0689_/S _0785_/S VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_143_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1065__C _1065_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_115_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1219_ VGND VPWR _1214_/X _1212_/X _1216_/X _1219_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_84_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1414__327 la_data_out[105] _1414__327/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_121_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_466 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_719 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input18_A la_data_in[49] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_29_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_835 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0616__A _0834_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_38_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_340 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_362 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_395 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_522 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1447__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_103_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_750 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0753__A1 _1102_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_67_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1004_ _1062_/D _1038_/D _1077_/B _1004_/D _1013_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_207_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_890 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_709 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0719_ _0746_/A _0742_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_1_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1092__A _1094_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_58_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1060 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1071 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_170 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_875 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0726__A1 _1057_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_82_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1484_ VGND VPWR _1484_/X _1484_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_140_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1151__A1 wb_clk_i VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_82_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_747 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_539 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input85_A wbs_dat_i[21] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_333 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_594 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1460__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1725 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_473 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0804__A _1497_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0984_ _0984_/Y _0984_/B _0984_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_164_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1467_ VGND VPWR _1467_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_476 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_837 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_358 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0626__A0 _1504_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_76_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1051__B1 _0848_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_155_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1455__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0965__A1_N _0869_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_135_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1321_ _1321_/Q _1253_/Y _1321_/D _1326_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_25_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1252_ VGND VPWR _1247_/X _1246_/X _1248_/X _1252_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XANTENNA__1106__A1 _1100_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1106__B2 _1065_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_209_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1183_ VGND VPWR _1180_/X _1179_/X _1181_/X _1183_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_64_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1715 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0865__B1 _0864_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_65_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_936 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0967_ _1141_/A _0997_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_140_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0898_ input90/X _0897_/X _0907_/A _0842_/X _0898_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_173_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput210 VPWR VGND la_data_out[9] _1483_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput221 VPWR VGND wbs_dat_o[18] _0688_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_66_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput232 VPWR VGND wbs_dat_o[28] _0635_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_86_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput243 VPWR VGND wbs_dat_o[9] _0735_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_153_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1341__254 la_data_out[32] _1341__254/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_183_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input48_A la_oenb[45] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0619__A _1021_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_93_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_741 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0821_ _0821_/B _0822_/D _0821_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_122_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1024__B1 _1010_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_116_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0752_ VGND VPWR _0752_/X _0752_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0801__B _1488_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0683_ VGND VPWR _0683_/X _0683_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1304_ _1304_/Q _1227_/Y _1304_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_211_1401 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1235_ VGND VPWR _1231_/X _1230_/X _1232_/X _1235_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_133_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1166_ VGND VPWR _1160_/X _1158_/X _1162_/X _1166_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_65_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1097_ _1481_/A _1097_/Y _1097_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_59_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1267__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_146_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_265 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input102_A wbs_dat_i[8] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_38_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1006__B1 _1005_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_50_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0902__A _0949_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_269 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_442 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output154_A _1490_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1020_ _1019_/Y _1015_/Y _1013_/Y _0832_/X _1018_/Y _1281_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41oi_4
XFILLER_130_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0783__S _1034_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0804_ _1495_/A _1496_/A _0805_/B _1494_/A _1497_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_50_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_781 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0735_ VGND VPWR _0735_/X _0735_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0666_ VGND VPWR _0666_/X _0666_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1218_ VGND VPWR _1214_/X _1212_/X _1216_/X _1218_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_168_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1149_ input72/X _1149_/X _1134_/B _0811_/A _1148_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_368 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0722__A _1485_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_120_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_935 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_946 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1347__260 la_data_out[38] _1347__260/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XANTENNA__0616__B _0834_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_204_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_330 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_341 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_352 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_396 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_272 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1463__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_140_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1003_ _1003_/Y _1003_/A _1003_/C _1003_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_110_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0807__A _1501_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_34_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1396__309 la_data_out[87] _1396__309/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_163_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1305__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_11_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0718_ VGND VPWR _0718_/X _0718_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0649_ VGND VPWR _0663_/S _0884_/A _1325_/Q _0650_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1083 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0680__A1 _0950_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0983__A2 _0824_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_120_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input30_A la_data_in[61] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_209_517 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_644 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_187 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1328__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_105_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_821 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_182 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1458__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_145_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_887 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0974__A2 _0824_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_103_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1483_ VGND VPWR _1483_/X _1483_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input78_A wbs_dat_i[15] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_551 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_325 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1908 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0983_ _0982_/X _0824_/X _0981_/Y _0990_/D input19/X _0984_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41oi_4
XANTENNA__0804__B _1496_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_203_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1188__A _1204_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_146_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1466_ VGND VPWR _1466_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_141_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1051__A1 _1026_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1320_ _1320_/Q _1252_/Y _1320_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_29_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1251_ VGND VPWR _1247_/X _1246_/X _1248_/X _1251_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_96_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1471__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1182_ VGND VPWR _1180_/X _1179_/X _1181_/X _1182_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_209_155 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1727 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_948 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0966_ _0966_/X _1097_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_203_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0897_ VGND VPWR _0897_/B _0897_/X _0820_/C _0897_/C VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_31_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput200 VPWR VGND la_data_out[29] _1503_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput211 VPWR VGND wbs_ack_o _1298_/Q VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput222 VPWR VGND wbs_dat_o[19] _0683_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_133_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput233 VPWR VGND wbs_dat_o[29] _0631_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_192_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1449_ VGND VPWR _1449_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_753 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1380__293 la_data_out[71] _1380__293/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_201_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_624 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0820_ _0820_/C _0906_/A _0821_/B _0820_/D _0820_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_200_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1024__A1 _1030_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_70_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0751_ VGND VPWR _0770_/S _1305_/Q _1102_/A _0752_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__1466__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_122_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0682_ VGND VPWR _0692_/S _1318_/Q _1493_/A _0683_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__0783__A0 _1140_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_171_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0801__C _1487_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_170_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1303_ _1303_/Q _1226_/Y _1303_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_57_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1234_ VGND VPWR _1231_/X _1230_/X _1232_/X _1234_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_49_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1165_ VGND VPWR _1160_/X _1158_/X _1162_/X _1165_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_64_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1096_ _1096_/Y _1096_/A _1143_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_20_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1364__277 la_data_out[55] _1364__277/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_139_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1397 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0949_ VPWR VGND _0949_/A _0999_/B VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_649 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_727 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0765__A0 _1477_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_50_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_944 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input60_A la_oenb[57] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output147_A _1474_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_182_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0803_ _1491_/A _1492_/A _0805_/A _1490_/A _1493_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XANTENNA__1196__A _1204_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_116_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0734_ VGND VPWR _0744_/S _1308_/Q _1059_/B _0735_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__0756__A0 _1109_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_115_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0665_ VGND VPWR _0665_/S _1321_/Q _1496_/A _0666_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_131_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1254 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1217_ _1216_/X _1217_/Y _1214_/X _1212_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_66_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_826 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1310 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1148_ _1148_/Y input1/X _0917_/B _0917_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1079_ _1082_/B _1079_/B _1079_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_59_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_counter.clk clkbuf_3_1_0_counter.clk/A _1322_/CLK VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_135_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_320 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_342 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_353 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_375 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_397 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1002_ _1034_/D _1002_/C _1073_/B _1003_/C _0817_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_2
XANTENNA__0807__B _1500_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_34_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0729__A0 _1067_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_102_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0717_ VGND VPWR _0717_/S _1311_/Q _1486_/A _0718_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_171_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0648_ VGND VPWR _0648_/X _0648_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_106_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_689 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0733__A _1483_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1420__333 la_data_out[111] _1420__333/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_167_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_711 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_722 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput100 VPWR VGND _1099_/A1 wbs_dat_i[6] VGND VPWR sky130_fd_sc_hd__buf_2
XANTENNA__1145__B1 _1140_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_799 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input23_A la_data_in[54] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_56_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_851 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_172 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__B1 _0958_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_560 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1474__A _1474_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1482_ VGND VPWR _1482_/X _1482_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_140_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1404__317 la_data_out[95] _1404__317/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_108_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0728__A _1484_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_58_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_147 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_118 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0638__A _1501_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_37_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1705 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1469__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0982_ _0982_/A _0982_/B _1092_/B _0982_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_18_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0804__C _1495_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_9_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1465_ VGND VPWR _1465_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1318__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_8_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_445 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input90_A wbs_dat_i[26] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_168_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output177_A _1482_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_170_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1250_ VGND VPWR _1247_/X _1246_/X _1248_/X _1250_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_1_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1181_ VPWR VGND _1205_/A _1181_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0865__A2 input93/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_64_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0965_ _1286_/D _0869_/X _0963_/Y _0964_/Y _0962_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_186_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0896_ VGND VPWR _0831_/Y _0889_/Y _1067_/A _0896_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_31_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput201 VPWR VGND la_data_out[2] _1476_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_192_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput212 VPWR VGND wbs_dat_o[0] _0784_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_173_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput223 VPWR VGND wbs_dat_o[1] _0778_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput234 VPWR VGND wbs_dat_o[2] _0771_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1448_ VGND VPWR _1448_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_114_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_526 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0856__A2 input95/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_83_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_916 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_408 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_960 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_146 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_537 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_920 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0651__A _1499_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_128_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0750_ _1047_/A _0770_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__1024__A2 _1050_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_200_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_953 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0681_ VGND VPWR _1319_/D _0681_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_155_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0801__D _1482_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_87_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1482__A _1482_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1302_ _1302_/Q _1225_/Y _1302_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_96_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1425 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1233_ VGND VPWR _1231_/X _1230_/X _1232_/X _1233_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_96_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1164_ VGND VPWR _1160_/X _1158_/X _1162_/X _1164_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_65_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0826__A _0834_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_25_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1095_ _1134_/B _1143_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_18_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1107__A2_N _1102_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_178_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0948_ _1142_/D _0948_/C _1142_/B _0948_/Y _0816_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_118_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0879_ _0907_/A _0879_/B _0958_/C _0879_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_134_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1006__A2 _1013_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_956 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input53_A la_oenb[50] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_84_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0646__A _1021_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1477__A _1477_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_0802_ _0949_/A _1038_/D _1004_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_204_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_790 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0733_ _1059_/B _1483_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_171_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0664_ VGND VPWR _1322_/D _0664_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_170_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1331__244 io_oeb[37] _1331__244/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_211_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1216_ VPWR VGND _1248_/A _1216_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1147_ _1267_/D _1027_/X _1144_/Y _1146_/Y _1140_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_25_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1322 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0692__A0 _0986_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1078_ _1078_/B _1078_/C _1077_/X _1082_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3b_1
XFILLER_74_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0747__A1 _1481_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_119_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_643 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_321 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_332 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_354 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_376 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_387 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_731 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1001_ _1001_/A _1094_/C _1001_/C _1094_/A _1003_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_47_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0807__C _1499_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_63_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1000__A _1111_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_163_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0716_ VGND VPWR _1312_/D _0716_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_132_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0647_ VGND VPWR _0665_/S _1325_/Q _0884_/A _0648_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_154_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0665__A0 _1496_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_657 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_896 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_395 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1145__A1 _1094_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xinput101 wbs_dat_i[7] _1096_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_118_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input16_A la_data_in[47] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_45_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_162 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_173 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1481_ VGND VPWR _1481_/X _1481_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1490__A _1490_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_94_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0895__B1 _0790_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0647__A0 _0884_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_165_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0834__A _0834_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_56_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_739 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1337__250 io_out[37] _1337__250/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_132_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input8_A la_data_in[39] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_98_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1063__B1 _1067_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0919__A _1080_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_209_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_498 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0981_ _0981_/A _0981_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_14_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0804__D _1494_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_146_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1485__A _1485_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_51_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_391 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1464_ VGND VPWR _1464_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0829__A _0841_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_25_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_829 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1066 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input83_A wbs_dat_i[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_128_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_102 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1180_ VPWR VGND _1204_/A _1180_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0964_ _0790_/A _0971_/D _0940_/C _0964_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_18_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0895_ _1293_/D _0887_/Y _0891_/A _0894_/Y _0790_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_146_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput202 VPWR VGND la_data_out[30] _1504_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_133_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput213 VPWR VGND wbs_dat_o[10] _0730_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_192_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput224 VPWR VGND wbs_dat_o[20] _0679_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_173_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput235 VPWR VGND wbs_dat_o[30] _0627_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_86_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1447_ VGND VPWR _1447_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_972 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_736 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_932 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1024__A3 _1050_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_196_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0680_ VGND VPWR _0689_/S _0950_/A _1319_/Q _0681_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_183_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1301_ _1301_/Q _1221_/Y _1301_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1232_ VGND VPWR _1232_/X _1248_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1163_ VGND VPWR _1160_/X _1158_/X _1162_/X _1163_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_93_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1094_ _1094_/B _1134_/B _1094_/A _1094_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_64_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1537 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0842__A _0945_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1308__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_197_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0947_ VPWR VGND _1142_/D _0947_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_147_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0878_ VPWR VGND _0958_/C _0945_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_173_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_401 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_968 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input46_A la_oenb[43] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0927__A _0938_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_46_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_552 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0801_ _1489_/A _1482_/A _1487_/A _1488_/A _1004_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_200_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0732_ VGND VPWR _1309_/D _0732_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_155_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0663_ VGND VPWR _0663_/S _1497_/A _1322_/Q _0664_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_115_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1493__A _1493_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_83_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1370__283 la_data_out[61] _1370__283/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_6_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1215_ VPWR VGND _1248_/A _1256_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_211_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0837__A _0891_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_65_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1146_ _0790_/A _1145_/Y _0980_/A _1146_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_1_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_327 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1334 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1077_ _1077_/A _1077_/X _1077_/B _1085_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_41_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_300 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input100_A wbs_dat_i[6] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_311 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_322 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_883 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_333 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_344 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_355 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_366 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1093__D1 _0997_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_199_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_377 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_388 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_399 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_743 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output152_A _1488_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_105_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1354__267 la_data_out[45] _1354__267/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_121_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1000_ _1003_/A _1111_/A _1000_/C _1000_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_47_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0807__D _1498_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1488__A _1488_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_76_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0715_ VGND VPWR _0715_/S _1030_/A _1312_/Q _0716_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_171_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0646_ VPWR VGND _0665_/S _1021_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_63_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1129_ _1129_/Y _1129_/A _1129_/C _1129_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_81_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput102 VPWR VGND _1079_/A wbs_dat_i[8] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_46_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_190 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1101__A _1118_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_38_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__A2 _1142_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_174 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_185 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_196 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1480_ VGND VPWR _1480_/X _1480_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0834__B _0834_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_165_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0629_ VGND VPWR _1329_/D _0629_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1063__A1 _1059_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_50_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_823 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0760__A _1478_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_202_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1138__A1_N _1027_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_120_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0935__A _1496_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_45_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0980_ _1000_/B _0980_/B _0984_/A _0980_/D _0980_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_53_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0670__A _1495_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_185_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0977__A1_N _0966_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1463_ VGND VPWR _1463_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1410__323 la_data_out[101] _1410__323/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_94_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_537 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0755__A _1479_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_2_1078 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_counter.clk clkbuf_2_3_0_counter.clk/A clkbuf_3_5_0_counter.clk/A VGND
+ VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0921__C _0921_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_182_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input76_A wbs_dat_i[13] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1559 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0963_ _0963_/Y _0963_/B _0963_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XANTENNA__1496__A _1496_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0894_ VGND VPWR _0894_/Y _0893_/X _0889_/Y _0849_/A _0891_/Y VGND VPWR sky130_fd_sc_hd__a31oi_1
XFILLER_185_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput203 VPWR VGND la_data_out[31] _1505_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput214 VPWR VGND wbs_dat_o[11] _0725_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_12_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput225 VPWR VGND wbs_dat_o[21] _0674_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_173_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput236 VPWR VGND wbs_dat_o[31] _0621_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1446_ VGND VPWR _1446_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_141_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_745 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_907 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_277 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0777__A0 _1132_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_139_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_550 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_200 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_748 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0932__B _0947_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_944 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1300_ _1300_/Q _1220_/Y _1300_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_65_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1231_ VPWR VGND _1247_/A _1231_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_211_1416 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1162_ VPWR VGND _1162_/A _1162_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1093_ _1118_/B _1085_/D _1091_/X _1108_/A _0997_/A _1093_/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_1516 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1549 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1345 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1003__B _1003_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_90_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1389 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0946_ _0993_/B _1000_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_146_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0877_ _0990_/D _0877_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_146_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_564 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_925 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input39_A la_oenb[36] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0927__B _0949_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_208_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_597 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0800_ _1486_/A _1483_/A _1484_/A _1485_/A _1038_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_204_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0731_ VGND VPWR _0742_/S _1067_/B _1309_/Q _0732_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_183_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0662_ VGND VPWR _0662_/X _0662_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1214_ _1247_/A _1214_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__0837__B _0884_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_38_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_807 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_818 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1145_ _1094_/B _1140_/B _1145_/Y _0842_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_20_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1076_ _1275_/D _1041_/X _1074_/Y _1070_/B _1075_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_20_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0929_ _0940_/C _0929_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_107_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_312 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_345 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_523 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_356 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_378 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0938__A _0938_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_67_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0714_ VGND VPWR _0714_/X _0714_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_171_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0645_ _0884_/A _1500_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_154_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1009__A _1486_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_615 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1128_ _1142_/D input4/X _1135_/B _1129_/C _0811_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_25_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1059_ _1059_/Y _1059_/B _1067_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_41_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_736 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput103 VPWR VGND _1072_/A wbs_dat_i[9] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_133_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_131 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_142 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_153 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_164 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_876 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1499__A _1499_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_719 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0834__C _0834_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_143_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0628_ VGND VPWR _0636_/S _1504_/A _1329_/Q _0629_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_63_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_106 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_835 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input21_A la_data_in[52] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_190_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1112__A _1112_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_53_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0951__A _0951_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_34_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1462_ VGND VPWR _1462_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1392__305 la_data_out[83] _1392__305/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_182_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input69_A la_oenb[66] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_194_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1433__346 la_data_out[124] _1433__346/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_137_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1709 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0962_ _0993_/B _0962_/B _0963_/B _0962_/D _0980_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_159_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0893_ input91/X _0892_/X _0918_/B _0842_/X _0893_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_88_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput204 VPWR VGND la_data_out[3] _1477_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput215 VPWR VGND wbs_dat_o[12] _0718_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_154_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput226 VPWR VGND wbs_dat_o[22] _0666_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput237 VPWR VGND wbs_dat_o[3] _0766_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_173_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1445_ VGND VPWR _1445_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0710__A1 _1010_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_55_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0701__A1 _0993_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_58_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output175_A _1480_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_136_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1230_ VPWR VGND _1246_/A _1230_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1161_ VPWR VGND _1256_/A _1162_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1092_ _1108_/A _1092_/B _1094_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_209_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_716 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0945_ _0993_/B _0982_/A _0945_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_186_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0876_ VPWR VGND _1142_/B _1080_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_106_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_716 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1891 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_165 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1266__RESET_B _1156_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_75_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_521 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_381 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1120__A _1120_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1398__311 la_data_out[89] _1398__311/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_106_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0730_ VGND VPWR _0730_/X _0730_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0661_ VGND VPWR _0665_/S _1322_/Q _1497_/A _0662_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_100_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_970 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1213_ VPWR VGND _1247_/A _1255_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0837__C _0888_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_93_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1144_ _1144_/Y _1144_/A _1144_/C _1144_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_1_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1075_ _1026_/A _1005_/X _1075_/Y _1062_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_209_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1358 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1030__A _1030_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_37_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0928_ _0945_/B _0877_/A _0982_/A _0824_/A _0940_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a22oi_4
XFILLER_146_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0859_ _1077_/B _1038_/D _0922_/A _1004_/D _1085_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_31_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1205__A _1205_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_79_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_830 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_302 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1870 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_324 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_346 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1297__D _1297_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_196_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input51_A la_oenb[48] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_175_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_550 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0713_ VGND VPWR _0717_/S _1312_/Q _1030_/A _0714_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_144_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0644_ VGND VPWR _1326_/D _0644_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1009__B _1485_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_83_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0898__B1 _0897_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_100_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1025__A _1050_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_2_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_605 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1099 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1127_ _1129_/B _1134_/B _1127_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_20_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1058_ _1057_/Y _1055_/Y _1054_/Y _0832_/X _1056_/Y _1277_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41oi_4
XFILLER_15_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_822 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1075__B1 _1005_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_179_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput104 VPWR VGND _1094_/B wbs_sel_i[0] VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_66_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0774__A _1475_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_44_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1066__B1 _0790_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_143 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_154 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_165 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_176 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_888 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input99_A wbs_dat_i[5] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__0959__A4 _1142_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_187 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_198 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1360__273 la_data_out[51] _1360__273/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_201_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0949__A _0949_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_84_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_181 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0627_ VGND VPWR _0627_/X _0627_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1344__257 la_data_out[35] _1344__257/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_50_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1063__A3 _1070_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_847 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0769__A _1476_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_172_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input14_A la_data_in[45] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_91_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1039__B1 _1005_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_92_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1461_ VGND VPWR _1461_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_114_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input6_A la_data_in[37] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_100_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1213__A _1255_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_82_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0962__A _0980_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0961_ VGND VPWR _0962_/B _0999_/B _1070_/A _0961_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_201_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_442 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0892_ VGND VPWR _0897_/B _0892_/X _0820_/D _0892_/C VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_185_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput205 VPWR VGND la_data_out[4] _1478_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_57_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput216 VPWR VGND wbs_dat_o[13] _0714_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput227 VPWR VGND wbs_dat_o[23] _0662_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_154_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput238 VPWR VGND wbs_dat_o[4] _0762_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_153_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1444_ VGND VPWR _1444_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1033__A _1033_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_64_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_725 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_358 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1283__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_23_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_881 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input81_A wbs_dat_i[18] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1400__313 la_data_out[91] _1400__313/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_196_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output168_A _1503_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_9_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1118__A _1118_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_65_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1160_ VPWR VGND _1160_/A _1160_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1091_ _1110_/A _1481_/A _1102_/A _1090_/X _1091_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_4_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_780 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0944_ _0944_/A _0944_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_72_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0875_ _1080_/A _0875_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_88_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0916__C1 _0980_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_115_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0695__A1 _0986_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_95_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1289_ _1497_/A _1200_/Y _1289_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_71_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_728 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_216 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_916 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0660_ VGND VPWR _1323_/D _0660_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_982 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1212_ VPWR VGND _1246_/A _1212_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1143_ _1144_/C _1143_/B _1143_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_38_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1074_ _1074_/Y _1074_/A _1074_/C _1074_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_93_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1348 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0927_ _0927_/X _0927_/C _0938_/A _0949_/A _0961_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_159_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0858_ _1085_/D _1062_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_162_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0789_ VPWR VGND _0790_/A _0861_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_115_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0668__A1 _1496_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_56_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_303 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_314 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1882 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_325 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_336 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_347 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_369 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input44_A la_oenb[41] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_171_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0659__A1 _0914_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_75_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_864 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_591 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0712_ _1030_/A _1487_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_89_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0643_ VGND VPWR _0663_/S _0891_/A _1326_/Q _0644_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_100_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1009__C _1484_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1025__B _1050_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_38_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1126_ _1129_/A _1141_/A _1126_/C _1141_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_25_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0864__B _0897_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_202_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1057_ _1057_/B _1057_/Y _1097_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_41_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1075__A1 _1026_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_834 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_333 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput105 _1016_/B wbs_sel_i[1] VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_62_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1216__A _1248_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_44_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1066__A1 input73/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_25_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_122 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_155 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0790__A _0790_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_73_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_166 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_177 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_188 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output150_A _1486_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1126__A _1141_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_27_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0626_ VGND VPWR _0639_/S _1329_/Q _1504_/A _0627_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_154_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0740__A0 _1050_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_100_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1109_ _1109_/A _1110_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_81_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1383__296 la_data_out[74] _1383__296/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_42_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_859 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1039__A1 _1026_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1460_ VGND VPWR _1460_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_153_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_529 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_counter.clk clkbuf_3_5_0_counter.clk/A _1294_/CLK VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_128_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0713__A0 _1030_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_86_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_601 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1507 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_409 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0960_ VPWR VGND _1070_/A _0985_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_60_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0891_ _0891_/B _0891_/Y _0891_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_179_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput206 VPWR VGND la_data_out[5] _1479_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_182_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput217 VPWR VGND wbs_dat_o[14] _0709_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_127_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput228 VPWR VGND wbs_dat_o[24] _0658_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput239 VPWR VGND wbs_dat_o[5] _0757_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_153_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1443_ VGND VPWR _1443_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_269 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1224__A _1248_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_58_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input109_A wbs_we_i VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_893 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input74_A wbs_dat_i[11] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_182_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1408 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1134__A _1134_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_37_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1090_ VPWR VGND _1090_/X _1478_/A _1109_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_92_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_792 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0943_ _0940_/Y _0848_/X _0942_/Y _0935_/Y _1288_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__a22oi_1
XFILLER_202_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0874_ _0874_/A _0874_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_146_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1044__A _1070_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_95_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1288_ _1496_/A _1199_/Y _1288_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_186_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1423__336 la_data_out[114] _1423__336/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_71_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0793__A _1503_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_74_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_243 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0968__A _0979_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_151_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_994 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1205 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1211_ VPWR VGND _1246_/A hold2/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_46_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1142_ _1142_/D input2/X _1142_/B _1144_/B _0811_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_37_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1073_ _1121_/D _1073_/C _1073_/B _1074_/C _0814_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_53_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0926_ _0961_/C _1491_/A _1493_/A _0979_/A _1490_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_88_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0857_ _0851_/Y _0848_/X _0856_/Y _0795_/A _1296_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__a22oi_1
XFILLER_88_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0788_ _1027_/A _0861_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_115_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0878__A _0945_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_130_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_604 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1761 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1502__A _1502_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_304 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1894 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_348 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input37_A la_oenb[34] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_681 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0840__A_N _1505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_389 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0711_ VGND VPWR _1313_/D _0711_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_183_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0642_ VPWR VGND _0663_/S _0785_/S VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_100_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0698__A _1047_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_112_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1009__D _1483_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_152_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0898__A2 input90/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_170_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1125_ _1126_/C _1132_/B _1125_/A _1125_/B _1132_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_93_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1056_ _1056_/Y _1056_/A _1072_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_20_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_846 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0909_ _0909_/Y _0909_/B _0909_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_107_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput106 VPWR VGND _0982_/A wbs_sel_i[2] VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_153_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1013 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1388__301 la_data_out[79] _1388__301/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_57_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_445 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_629 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1232__A _1248_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1429__342 la_data_out[120] _1429__342/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_72_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_651 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_112 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1691 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_695 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_134 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_145 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_156 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_167 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1311__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__A1_N _0869_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_144_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0625_ VGND VPWR _1330_/D _0625_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1108_ _1108_/A _1141_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_54_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0891__A _0891_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1039_ _1026_/A _1005_/X _1039_/Y _1038_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_41_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0731__A1 _1067_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_88_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0976__A _1493_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_190_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_877 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_470 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1047__A _1047_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_144_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1350__263 la_data_out[41] _1350__263/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0796__A _1477_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_1_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0890_ _1500_/A _0891_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_35_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput207 VPWR VGND la_data_out[6] _1480_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_142_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_661 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput218 VPWR VGND wbs_dat_o[15] _0704_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_182_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput229 VPWR VGND wbs_dat_o[25] _0653_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_153_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0943__A1 _0848_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1442_ VGND VPWR _1442_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1334__247 io_out[34] _1334__247/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_4_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_327 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1505__A _1505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_82_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1240__A _1248_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input67_A la_oenb[64] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_151_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1509 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0973__B _0973_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_45_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0942_ _0942_/Y _1005_/A _1001_/A _0872_/B _0941_/X input86/X VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a311oi_4
XFILLER_53_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0873_ _0873_/C _1078_/C _0881_/A _0873_/D _0873_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_88_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_981 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1287_ _1495_/A _1198_/Y _1287_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_55_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1060__A _1477_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_63_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_557 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output173_A _1478_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_112_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0968__B _0986_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_151_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1210_ VGND VPWR _1204_/X _1203_/X _1205_/X _1210_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_113_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1141_ _1144_/A _1141_/A _1141_/C _1141_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_187_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1072_ _1074_/B _1072_/B _1072_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_207_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0925_ VGND VPWR _0927_/C _0951_/A _1496_/A _0950_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_120_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0856_ _0856_/Y _1005_/A _0918_/B _0872_/B _0855_/X input95/X VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a311oi_4
XFILLER_106_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0787_ VPWR VGND _0787_/A _1027_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1011__B1 _1489_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_115_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_316 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_338 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0710_ VGND VPWR _0715_/S _1010_/A _1313_/Q _0711_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0979__A _0979_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_0641_ _0746_/A _0785_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_143_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1124_ _1270_/D _1041_/X _1122_/Y _1115_/A _1123_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_54_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1055_ _0814_/D _1055_/Y _1055_/B _1065_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3b_4
XFILLER_53_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_858 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0908_ _0907_/X _0824_/X _0906_/Y _0990_/D input26/X _0909_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41oi_4
XFILLER_198_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0839_ _0889_/B _0873_/A _0839_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_200_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput107 VPWR VGND _0841_/A wbs_sel_i[3] VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_44_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1025 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1058 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_663 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1681 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_168 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_545 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_740 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1142__B _1142_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_188_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0624_ VGND VPWR _0636_/S _1505_/A _1330_/Q _0625_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1107_ _0832_/X _1272_/D VGND VPWR _1106_/Y _1099_/Y _1102_/A VGND VPWR sky130_fd_sc_hd__a2bb2oi_1
XFILLER_93_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1038_ _1085_/D _1062_/A _1038_/X _1118_/B _1038_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_22_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1286__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_210_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_405 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input97_A wbs_dat_i[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_160_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1153__A hold3/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_76_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0895__A2_N _0891_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_91_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_670 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1149__A1_N input72/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_199_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_669 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1238__A _1246_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_87_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1301__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_118_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0796__B _1476_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_89_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_389 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0988__A1_N _0966_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_725 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_736 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input12_A la_data_in[43] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_57_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput208 VPWR VGND la_data_out[7] _1481_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_126_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput219 VPWR VGND wbs_dat_o[16] _0700_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_142_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1441_ VGND VPWR _1441_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_142_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1373__286 la_data_out[64] _1373__286/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_190_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1061 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input4_A la_data_in[35] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_86_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_227 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_923 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0689__A1 _0979_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_89_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0941_ VGND VPWR _0947_/A _0941_/X _0816_/C _0941_/C VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_92_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0872_ _0873_/C _0872_/B _0918_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_35_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1900 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1922 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1286_ _1494_/A _1194_/Y _1286_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_186_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_461 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1840 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1129__C _1129_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_67_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output166_A _1501_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_97_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1140_ VPWR VGND _1141_/C _1140_/B _1140_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_37_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_66 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1071_ _1074_/A _1111_/A _1071_/C _1078_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_4_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1161__A _1256_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_207_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_580 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0924_ _1290_/D _0869_/X _0921_/Y _0915_/D _0923_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_14_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0855_ _0819_/C _0855_/X _0855_/C _0947_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_88_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1379__292 la_data_out[70] _1379__292/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_0786_ VGND VPWR _1299_/D _0786_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0770__A0 _1125_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_170_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1269_ _1477_/A _1165_/Y _1269_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1071__A _1111_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_45_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_306 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_328 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1246__A _1246_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_10_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0761__A0 _1118_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_823 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_878 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0640_ VGND VPWR _0640_/X _0640_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1156__A _1156_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_28_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1413__326 la_data_out[104] _1413__326/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_61_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1015 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1037 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1048 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1123_ _1100_/Y _0861_/X _1123_/Y _1118_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_93_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1054_ _1054_/C _1054_/B _1054_/Y _1054_/D _1078_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_39_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0907_ _0907_/B _0907_/X _0907_/A _0958_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_120_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0838_ _0985_/A _0914_/A _0889_/B _0838_/D _0949_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4_2
XFILLER_162_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0769_ VPWR VGND _1125_/B _1476_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_115_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput108 VPWR VGND _0834_/A wbs_stb_i VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_44_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_815 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_114 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_136 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_158 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0734__A0 _1059_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_133_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input42_A la_oenb[39] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_686 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_697 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0623_ _0636_/S _0746_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_98_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1150__B1 _1027_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1106_ _1105_/X _1100_/Y _1065_/C _1104_/X _1106_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22oi_1
XFILLER_54_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1037_ VPWR VGND _1118_/B _1077_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0964__B1 _0790_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_107_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput90 VPWR VGND input90/X wbs_dat_i[26] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_159_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_877 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_802 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1419__332 la_data_out[110] _1419__332/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_208_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1123__B1 _0861_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0796__C _1475_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1254__A hold2/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_172_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_748 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput209 VPWR VGND la_data_out[8] _1482_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_127_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1440_ VGND VPWR _1440_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_175_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_632 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0897__B _0897_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_8_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_935 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1299__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_202_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0940_ _0940_/B _0940_/C _0927_/X _0940_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3b_1
XFILLER_60_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0871_ VPWR VGND _1078_/C _0952_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_158_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1159__A _1255_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1340__253 irq[2] _1340__253/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_35_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0998__A _1490_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_66_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1285_ _1493_/A _1193_/Y _1285_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_68_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_440 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_732 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1069__A _1483_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_865 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input107_A wbs_sel_i[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_187_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_776 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input72_A wbs_dat_i[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_171_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1020__A2 _1015_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_97_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output159_A _1494_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_191_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1442__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1314__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1070_ VGND VPWR _1071_/C _1070_/B _1070_/A _1070_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_207_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_529 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0923_ _0849_/X _0910_/X _0923_/Y _0922_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_202_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0854_ VPWR VGND _0947_/A _0854_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_11_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0785_ VGND VPWR _0785_/S _1140_/B _1299_/Q _0786_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__1011__A2 _0938_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_143_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_counter.clk clkbuf_0_counter.clk/X clkbuf_2_3_0_counter.clk/A VGND VPWR
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_170_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1055__C _1065_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_170_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1268_ _1476_/A _1164_/Y _1268_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_186_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1199_ VGND VPWR _1196_/X _1195_/X _1197_/X _1199_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_129_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_307 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_318 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_518 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_76 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_835 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1437__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_119_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1027 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1172__A _1256_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_187_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1122_ _1122_/Y _1122_/A _1122_/C _1122_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_66_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1053_ VGND VPWR _1077_/A _0938_/A _1059_/B _1054_/D _1057_/B _1484_/A VGND VPWR
+ sky130_fd_sc_hd__a41o_1
XFILLER_4_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_304 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0906_ _0906_/A _0906_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_30_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0837_ _0839_/A _0891_/A _0888_/A _0884_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_179_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0768_ VGND VPWR _1302_/D _0768_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_130_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0699_ VGND VPWR _0717_/S _1315_/Q _0993_/D _0700_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_115_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput109 _0834_/C wbs_we_i VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_170_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_104 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_827 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_148 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1395__308 la_data_out[86] _1395__308/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_197_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1436__349 la_data_out[127] _1436__349/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_180_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_764 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input35_A la_oenb[32] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1142__D _1142_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0622_ _0834_/A _0746_/A _0787_/A _0834_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_98_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1150__B2 _1140_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_113_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1105_ VPWR VGND _1105_/X input7/X _0810_/C VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_38_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1036_ _1077_/A _1062_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_39_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_624 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0661__A0 _1497_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_22_657 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_808 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput80 VGND VPWR _0989_/A wbs_dat_i[17] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_174_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput91 wbs_dat_i[27] input91/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_122_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1391 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_counter.clk clkbuf_3_3_0_counter.clk/A _1326_/CLK VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0652__A0 _0888_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_9_617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_333 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_814 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1450__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_188_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_160 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1123__A1 _1100_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_187_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0882__B1 _0848_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_148_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_922 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1019_ _1489_/A _1019_/Y _1067_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_168_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0634__A0 _1502_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_168_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0796__D _1474_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_49_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0928__A1 _0982_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__0928__B2 _0877_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_126_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1445__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_141_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_644 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1180__A _1204_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_75_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1499_ VGND VPWR _1499_/X _1499_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1090__A _1109_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_27_535 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_914 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_947 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1099__B1 _0848_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_58_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0846__B1 _0790_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_79_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0870_ VGND VPWR _0917_/B _0917_/A _0824_/A _0952_/A VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_35_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1023__B1 _0824_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_31_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1284_ _1492_/A _1192_/Y _1284_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_42_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0999_ VGND VPWR _1000_/C _0999_/B _1050_/B _0999_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_10_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1266__CLK _1279_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_204_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1363__276 la_data_out[54] _1363__276/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_208_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_265 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input65_A la_oenb[62] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_486 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0922_ _0922_/Y _0922_/B _0922_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_140_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0853_ VPWR VGND _0872_/B _1092_/B VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_174_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0784_ VGND VPWR _0784_/X _0784_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput1 VGND VPWR input1/X la_data_in[32] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1267_ _1475_/A _1163_/Y _1267_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_84_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1289__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1198_ VGND VPWR _1196_/X _1195_/X _1197_/X _1198_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_37_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_308 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0712__A _1487_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0831__A2_N _0824_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_49_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0846__A2_N _1505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_87_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1147__A1_N _1027_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_210_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0622__A _0787_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_109_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output171_A _1505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_119_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1453__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_61_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1121_ _1121_/D input5/X _1135_/B _1122_/C _0810_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_43_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1052_ _1278_/D _1041_/X _1049_/Y _1051_/Y _1044_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_207_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_806 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0905_ _0980_/A _0903_/X _0828_/X _0830_/Y _0922_/B _0909_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_174_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0924__A1_N _0869_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0836_ _0945_/B _0877_/A _0841_/A _0824_/A _0849_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a22oi_4
XFILLER_190_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0767_ VGND VPWR _0767_/S _1477_/A _1302_/Q _0768_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_85_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0698_ VPWR VGND _0717_/S _1047_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_170_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1319_ _1319_/Q _1251_/Y _1319_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0707__A _1488_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_138 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1304__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput190 VPWR VGND la_data_out[1] _1475_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_43_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_776 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input28_A la_data_in[59] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_87_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1369__282 la_data_out[60] _1369__282/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_43_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_850 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_832 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1448__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_160_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0621_ VGND VPWR _0621_/X _0621_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_570 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1104_ _1104_/X _1118_/B _1103_/X _1115_/A _1102_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_19_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1035_ _1035_/Y _1035_/A _1035_/C _1035_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_35_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_636 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1327__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_206_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_680 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput70 wb_rst_i input70/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput81 wbs_dat_i[18] _0982_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_0819_ _0819_/C _0819_/B _0821_/A _0819_/D _0874_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_200_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput92 wbs_dat_i[28] _0879_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_89_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1403__316 la_data_out[94] _1403__316/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_41_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_573 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_826 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0643__A1 _0891_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1018_ _1018_/Y _1018_/A _1072_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_23_934 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input95_A wbs_dat_i[30] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0928__A2 _0945_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_181_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1461__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1053 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_948 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1074__C _1074_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_99_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1498_ VGND VPWR _1498_/X _1498_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1090__B _1478_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_64_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__B1 _0636_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_123_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1099__A1 _1099_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input10_A la_data_in[41] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_79_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1409__322 la_data_out[100] _1409__322/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1023__A1 _1016_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_196_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1023__B2 _1021_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1456__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_157_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1283_ _1491_/A _1191_/Y _1283_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_23_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0998_ _1490_/A _0999_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_14_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input2_A la_data_in[33] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_86_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_299 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1020__A4 _0832_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_163_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input58_A la_oenb[55] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_78_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_812 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1181 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0921_ _0921_/Y _0921_/A _0921_/C _0921_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_92_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0852_ _0852_/A _1092_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0783_ VGND VPWR _1034_/D _1299_/Q _1140_/B _0784_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_196_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1733 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput2 VGND VPWR input2/X la_data_in[33] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1266_ _1474_/A _1156_/A _1266_/D _1279_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_83_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_261 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1811 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1197_ VGND VPWR _1197_/X _1205_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_52_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1386__299 la_data_out[77] _1386__299/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_52_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1662 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1096__A _1096_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_69_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0903__A _0914_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_180_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0622__B _0834_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_158_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output164_A _1499_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_158_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1120_ _1122_/B _1143_/B _1120_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_43_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_631 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1051_ _1026_/A _0848_/X _1051_/Y _1054_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_59_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0904_ VPWR VGND _0980_/A _0952_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_50_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0835_ _0945_/B _0852_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0766_ VGND VPWR _0766_/X _0766_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0697_ VPWR VGND _0993_/D _1490_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_143_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1082__C _1082_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_61_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1318_ _1318_/Q _1250_/Y _1318_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_211_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0900__B1 _0790_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_22_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1563 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1249_ VGND VPWR _1247_/X _1246_/X _1248_/X _1249_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_38_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0723__A _1047_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_90_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput180 VPWR VGND la_data_out[10] _1484_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput191 VPWR VGND la_data_out[20] _1494_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_862 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_844 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_855 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0620_ VGND VPWR _0639_/S _1330_/Q _1505_/A _0621_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_109_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1279__CLK _1279_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_140_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1464__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_180_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1103_ _1090_/X _1110_/A _1480_/A _1103_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_187_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_472 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1034_ _1034_/D _1034_/C _1073_/B _1035_/C _0813_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_39_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1131__A1_N _1027_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_692 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput60 VGND VPWR _0906_/A la_oenb[57] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput71 VPWR VGND _0834_/B wbs_cyc_i VGND VPWR sky130_fd_sc_hd__buf_4
X_0818_ _0818_/B _0822_/C _0818_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
Xinput82 wbs_dat_i[19] _0973_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput93 wbs_dat_i[29] input93/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_85_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0749_ _1102_/A _1480_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_46_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_475 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input40_A la_oenb[37] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_164_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_585 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1459__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_203_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_681 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1017_ VPWR VGND _1079_/B _1072_/B VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
X_1426__339 la_data_out[117] _1426__339/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_39_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_946 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1088__B _1094_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input88_A wbs_dat_i[24] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_194_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_883 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1043 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1189__A _1205_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_189_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1497_ VGND VPWR _1497_/X _1497_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_113_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__A1 _0790_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_163_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_647 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1472__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_150_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1282_ _1490_/A _1190_/Y _1282_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_205_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1855 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_713 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0997_ _1111_/A _0997_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_101_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_290 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_389 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0920_ _1034_/D _0920_/C _1073_/B _0921_/C _0820_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_2
XFILLER_42_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0851_ _0809_/A _0809_/B _0851_/Y _0850_/Y _0849_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_1
XFILLER_31_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1467__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_122_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0782_ _1140_/B _1132_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_750 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1265_ VGND VPWR _1160_/A _1158_/A _1162_/A _1265_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_42_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput3 VGND VPWR input3/X la_data_in[34] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_84_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1196_ VPWR VGND _1204_/A _1196_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1834 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1674 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0994__A1 _0989_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_140_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0682__A0 _1493_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_input105_A wbs_sel_i[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_150_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0903__B _0938_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0622__C _0834_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input70_A wb_rst_i VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_158_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_720 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output157_A _1493_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_643 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1050_ _1054_/B _1050_/A _1050_/C _1050_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_130_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_131 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0673__A0 _0951_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_893 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0903_ _0903_/X _0992_/B _0914_/A _0938_/A _0903_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_119_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1197__A _1205_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_50_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0834_ VGND VPWR _0852_/A _0834_/B _0834_/A _0834_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_11_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0765_ VGND VPWR _0770_/S _1302_/Q _1477_/A _0766_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0696_ VGND VPWR _1316_/D _0696_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1353__266 la_data_out[44] _1353__266/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_9_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1317_ _1317_/Q _1249_/Y _1317_/D _1326_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1248_ VPWR VGND _1248_/A _1248_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_613 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1179_ VPWR VGND _1203_/A _1179_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1493 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput170 VPWR VGND io_out[30] _1504_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_122_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput181 VPWR VGND la_data_out[11] _1485_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput192 VPWR VGND la_data_out[21] _1495_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0914__A _0914_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_178_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_47 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1480__A _1480_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1102_ _1102_/Y _1109_/A _1102_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_81_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0808__B _0949_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_207_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1033_ _1035_/B _1072_/B _1033_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_35_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput50 VGND VPWR _0813_/D la_oenb[47] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput61 VGND VPWR _0820_/C la_oenb[58] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0817_ _0981_/A _0817_/B _0818_/B _0972_/A _0817_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_128_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput72 VPWR VGND input72/X wbs_dat_i[0] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_176_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput83 VPWR VGND _1143_/A wbs_dat_i[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xinput94 wbs_dat_i[2] _1134_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_137_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0748_ VGND VPWR _1306_/D _0748_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_107_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0679_ VGND VPWR _0679_/X _0679_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_130_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input33_A la_data_in[64] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_597 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_631 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1053__B1 _1057_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_12_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_686 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1475__A _1475_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_67_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_892 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1016_ VGND VPWR _1079_/B _1016_/B _1094_/A _1094_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_39_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_468 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1359__272 la_data_out[50] _1359__272/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_137_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1269__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_590 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1077 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1496_ VGND VPWR _1496_/X _1496_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_527 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_845 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0791__A2 _1298_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_159_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0922__A _0922_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_186_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1281_ _1489_/A _1186_/Y _1281_/D _1281_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_81_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1128 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1867 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_747 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0996_ _1283_/D _0966_/X _0994_/Y _0992_/C _0995_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_140_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_781 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_280 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1479_ VGND VPWR _1479_/X _1479_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_530 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1307__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_563 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0850_ _0850_/Y _0873_/D _0795_/B _0809_/B _0795_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
XFILLER_70_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0781_ VGND VPWR _1132_/C _1474_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1483__A _1483_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1264_ VGND VPWR _1160_/A _1158_/A _1162_/A _1264_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_83_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput4 VGND VPWR input4/X la_data_in[35] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0827__A _0834_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_36_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1195_ VPWR VGND _1203_/A _1195_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1824 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_566 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0979_ _0979_/A _0980_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_69_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input63_A la_oenb[60] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1478__A _1478_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_147_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0902_ _0949_/A _0992_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0833_ VGND VPWR _0831_/Y _0809_/Y _0832_/X _0833_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_50_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0764_ VGND VPWR _1303_/D _0764_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0695_ VGND VPWR _0715_/S _0986_/A _1316_/Q _0696_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_157_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1316_ _1316_/Q _1245_/Y _1316_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_9_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1247_ VPWR VGND _1247_/A _1247_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1178_ VGND VPWR _1171_/X _1169_/X _1173_/X _1178_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_37_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1632 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput160 VPWR VGND io_out[21] _1495_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_161_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput171 VPWR VGND io_out[31] _1505_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput182 VPWR VGND la_data_out[12] _1486_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_121_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput193 VPWR VGND la_data_out[22] _1496_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_135 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1376__289 la_data_out[67] _1376__289/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_124_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1101_ _1118_/A _1115_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_130_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1032_ _1035_/A _1111_/A _1032_/C _1078_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_207_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_190 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput40 VGND VPWR _0810_/B la_oenb[37] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_174_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0816_ _0816_/C _0816_/B _0818_/A _0816_/D _0957_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_190_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput51 VGND VPWR _0817_/A la_oenb[48] VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput62 VGND VPWR _0820_/D la_oenb[59] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput73 VPWR VGND input73/X wbs_dat_i[10] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_50_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput84 wbs_dat_i[20] _0958_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_89_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput95 VPWR VGND input95/X wbs_dat_i[30] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_190_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0747_ VGND VPWR _0767_/S _1481_/A _1306_/Q _0748_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_137_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0678_ VGND VPWR _0692_/S _1319_/Q _0950_/A _0679_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_118_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0750__A _1047_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0909__B _0909_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_input26_A la_data_in[57] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_87_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0628__A1 _1504_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__0925__A _1496_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_75_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1053__A1 _1484_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_156_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1491__A _1491_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0867__B2 _0790_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_67_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1015_ _0813_/D _1015_/Y _1015_/B _1065_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3b_4
XFILLER_35_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_852 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_863 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1067 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_280 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_291 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1486__A _1486_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_200_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1391__304 la_data_out[82] _1391__304/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_67_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1495_ VGND VPWR _1495_/X _1495_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_141_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1432__345 la_data_out[123] _1432__345/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_80_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input93_A wbs_dat_i[29] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_977 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1416__329 la_data_out[107] _1416__329/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_68_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1280_ _1488_/A _1185_/Y _1280_/D _1281_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_95_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1879 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0995_ _0929_/X _0910_/X _0995_/Y _0970_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_160_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1478_ VGND VPWR _1478_/X _1478_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_804 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_687 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_958 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_837 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0780_ VGND VPWR _1300_/D _0780_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_763 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1263_ VGND VPWR _1160_/A _1158_/A _1162_/A _1263_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_133_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput5 VGND VPWR input5/X la_data_in[36] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_65_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1194_ VGND VPWR _1188_/X _1187_/X _1189_/X _1194_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_149_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1858 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1397__310 la_data_out[88] _1397__310/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_578 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0978_ _0980_/B _0992_/A _0986_/A _1490_/A _0992_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_9_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_538 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input56_A la_oenb[53] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_78_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0901_ _0938_/A _0901_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_147_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0832_ VPWR VGND _0832_/X _1027_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_50_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0763_ VGND VPWR _0767_/S _1118_/A _1303_/Q _0764_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1494__A _1494_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_116_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_582 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0694_ VPWR VGND _0715_/S _0746_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_142_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0838__A _0914_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1315_ _1315_/Q _1244_/Y _1315_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_57_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1246_ VPWR VGND _1246_/A _1246_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1177_ VGND VPWR _1171_/X _1169_/X _1173_/X _1177_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_52_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1644 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_832 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1154__A_N input70/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput150 VPWR VGND io_out[12] _1486_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_118_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput161 VPWR VGND io_out[22] _1496_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_121_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput172 VPWR VGND io_out[3] _1477_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_161_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput183 VPWR VGND la_data_out[13] _1487_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput194 VPWR VGND la_data_out[23] _1497_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_153_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_158 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output162_A _1497_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1100_ _0958_/C _0947_/A _1094_/B _1080_/A _1100_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a22oi_4
XFILLER_43_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1031_ _1032_/C _1070_/C _1070_/A _1031_/B _1031_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_59_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1489__A _1489_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_146_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1001__B _1094_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_50_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput30 VGND VPWR _0864_/C la_data_in[61] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0840__B _1504_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xinput41 VGND VPWR _0810_/C la_oenb[38] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0815_ _0815_/B _0822_/B _0815_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_50_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput52 VGND VPWR _0817_/B la_oenb[49] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_174_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput63 VGND VPWR _0874_/A la_oenb[60] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_190_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput74 VPWR VGND _1056_/A wbs_dat_i[11] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_102_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput85 VGND VPWR _0944_/A wbs_dat_i[21] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0746_ VPWR VGND _0767_/S _0746_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xinput96 wbs_dat_i[31] input96/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_66_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0677_ VPWR VGND _0950_/A _1494_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_143_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1229_ VGND VPWR _1223_/X _1222_/X _1224_/X _1229_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_84_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_806 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_828 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input19_A la_data_in[50] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_63_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_445 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0925__B _0951_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1102__A _1102_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1343__256 la_data_out[34] _1343__256/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_8_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1053__A2 _1059_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1014_ _0917_/A _0917_/B _0824_/A _1065_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_207_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1012__A _1016_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_206_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0729_ VGND VPWR _0744_/S _1309_/Q _1067_/B _0730_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_669 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_875 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0936__A _0951_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_743 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0671__A _0897_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_292 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0785__A1 _1140_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_103_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1494_ VGND VPWR _1494_/X _1494_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input86_A wbs_dat_i[22] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0767__A1 _1477_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_103_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1330__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_64_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1349__262 la_data_out[40] _1349__262/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_79_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1497__A _1497_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_203_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0994_ _0989_/Y _1000_/B _0994_/Y _0993_/Y _0990_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_1
XFILLER_164_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0758__A1 _1109_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_30_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1477_ VGND VPWR _1477_/X _1477_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0930__A1 _1497_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_80_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_counter.clk clkbuf_3_7_0_counter.clk/A _1281_/CLK VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_83_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_775 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1262_ VGND VPWR _1160_/A _1158_/A _1162_/A _1262_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_211_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput6 VGND VPWR input6/X la_data_in[37] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_49_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1193_ VGND VPWR _1188_/X _1187_/X _1189_/X _1193_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_64_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_860 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_381 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0843__B _0877_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0977_ _1285_/D _0966_/X _0975_/Y _0964_/Y _0976_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_9_580 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_863 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_557 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1147__B2 _1146_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_78_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input49_A la_oenb[46] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0900_ _1292_/D _0896_/Y _0884_/A _0899_/Y _0790_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_37_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0831_ _0830_/Y _0831_/Y _1021_/B _0824_/X _0828_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_2
XFILLER_31_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0762_ VGND VPWR _0762_/X _0762_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0693_ VGND VPWR _0693_/X _0693_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1314_ _1314_/Q _1243_/Y _1314_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_111_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1245_ VGND VPWR _1239_/X _1238_/X _1240_/X _1245_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_2_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1176_ VGND VPWR _1171_/X _1169_/X _1173_/X _1176_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_65_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1656 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput140 VPWR VGND io_oeb[3] _1440_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput151 VPWR VGND io_out[13] _1487_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput162 VPWR VGND io_out[23] _1497_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_118_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput173 VPWR VGND io_out[4] _1478_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_121_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput184 VPWR VGND la_data_out[14] _1488_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput195 VPWR VGND la_data_out[24] _1498_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input103_A wbs_dat_i[9] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_71_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output155_A _1491_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_78_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1030_ _1030_/A _1031_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_130_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1001__C _1001_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_148_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput20 VGND VPWR input20/X la_data_in[51] VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput31 VGND VPWR _0855_/C la_data_in[62] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0814_ _0814_/C _0814_/B _0815_/B _0814_/D _0814_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XANTENNA__0840__C _1503_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xinput42 VGND VPWR _1088_/A la_oenb[39] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput53 VGND VPWR _0981_/A la_oenb[50] VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput64 VGND VPWR _0819_/B la_oenb[61] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_174_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput75 wbs_dat_i[12] _1046_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_196_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput86 input86/X wbs_dat_i[22] VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_0745_ VGND VPWR _0745_/X _0745_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_171_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput97 wbs_dat_i[3] _1127_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_176_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0676_ VGND VPWR _1320_/D _0676_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1228_ VGND VPWR _1223_/X _1222_/X _1224_/X _1228_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_113_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1159_ VPWR VGND _1255_/A _1160_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1453 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0925__C _0950_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_71_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1102__B _1109_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_38_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1382__295 la_data_out[73] _1382__295/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_169_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0941__B _0947_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_185_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_678 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_884 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1013_ _1013_/B _1078_/C _1013_/Y _1054_/C _1013_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4_2
XFILLER_81_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0728_ _1067_/B _1484_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_89_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0659_ VGND VPWR _0663_/S _0914_/A _1323_/Q _0660_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_98_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1203__A _1203_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_148_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1366__279 la_data_out[57] _1366__279/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_144_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input31_A la_data_in[62] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_209_617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_755 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_271 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_282 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_692 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1493_ VGND VPWR _1493_/X _1493_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0942__C1 _0941_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_141_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_837 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0933__C1 _0932_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_8_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_257 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1282__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_210_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input79_A wbs_dat_i[16] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_662 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0947__A _0947_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_739 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0993_ _0993_/C _0993_/B _0993_/Y _0993_/D _0997_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_203_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_counter.clk clkbuf_2_1_0_counter.clk/A clkbuf_3_3_0_counter.clk/A VGND
+ VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1018__A _1018_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_119_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1476_ VGND VPWR _1476_/X _1476_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_992 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1422__335 la_data_out[113] _1422__335/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_41_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_750 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_787 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1330_ _1330_/Q _1265_/Y _1330_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_123_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1261_ VGND VPWR _1255_/X _1254_/X _1256_/X _1261_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XANTENNA__0677__A _1494_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_96_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput7 VGND VPWR input7/X la_data_in[38] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1192_ VGND VPWR _1188_/X _1187_/X _1189_/X _1192_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_49_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1849 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0976_ _1493_/A _0976_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_118_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1459_ VGND VPWR _1459_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1406__319 la_data_out[97] _1406__319/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_19_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1211__A hold2/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_58_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1320__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_191_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0830_ _0907_/A _0830_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_70_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0761_ VGND VPWR _0770_/S _1303_/Q _1118_/A _0762_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_155_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0692_ VGND VPWR _0692_/S _1316_/Q _0986_/A _0693_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_170_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1313_ _1313_/Q _1242_/Y _1313_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_110_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1513 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0838__C _0949_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1244_ VGND VPWR _1239_/X _1238_/X _1240_/X _1244_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_133_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0649__A1 _0884_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_49_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1175_ VGND VPWR _1171_/X _1169_/X _1173_/X _1175_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_20_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1668 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1442 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1031__A _1070_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_107_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0959_ _0958_/X _1142_/B _0957_/Y _1142_/D input21/X _0963_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41oi_4
XFILLER_119_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput130 VPWR VGND io_oeb[28] _1465_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_118_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput141 VPWR VGND io_oeb[4] _1441_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput152 VPWR VGND io_out[14] _1488_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_157_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_705 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput163 VPWR VGND io_out[24] _1498_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput174 VPWR VGND io_out[5] _1479_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_716 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput185 VPWR VGND la_data_out[15] _1489_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput196 VPWR VGND la_data_out[25] _1499_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input61_A la_oenb[58] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_194_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output148_A _1484_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_79_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1387__300 la_data_out[78] _1387__300/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_143_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1089 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1428__341 la_data_out[119] _1428__341/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_146_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1001__D _1094_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_147_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput10 VGND VPWR _1073_/C la_data_in[41] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_163_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput21 VGND VPWR input21/X la_data_in[52] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0813_ _0813_/C _0813_/B _0815_/A _0813_/D _0813_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_141_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput32 VGND VPWR _0843_/C la_data_in[63] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_156_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput43 VGND VPWR _0814_/A la_oenb[40] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0840__D _1502_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xinput54 VGND VPWR _0972_/A la_oenb[51] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput65 VGND VPWR _0819_/C la_oenb[62] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0744_ VGND VPWR _0744_/S _1306_/Q _1481_/A _0745_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput76 wbs_dat_i[13] _1033_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_157_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_893 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xinput87 input87/X wbs_dat_i[23] VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput98 VPWR VGND _1120_/A wbs_dat_i[4] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_171_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_392 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0675_ VGND VPWR _0689_/S _0951_/A _1320_/Q _0676_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_66_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1026__A _1026_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_57_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1227_ VGND VPWR _1223_/X _1222_/X _1224_/X _1227_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_42_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1158_ VPWR VGND _1158_/A _1158_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1432 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1465 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1089_ _1110_/A _1475_/A _1477_/A _1476_/A _1474_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_59_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_557 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_753 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_420 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_624 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1053__A4 _0938_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_129_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1012_ _1054_/C _1092_/B _1016_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_130_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_285 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0624__S _0636_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_148_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0727_ VGND VPWR _1310_/D _0727_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0658_ VGND VPWR _0658_/X _0658_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0996__A1_N _0966_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_27_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1251 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0934__A1_N _0832_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_167_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_126 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_387 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0703__A0 _1489_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_76_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input24_A la_data_in[55] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_250 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_283 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_294 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1492_ VGND VPWR _1492_/X _1492_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_140_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0933__B1 _0790_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_137_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1333__246 io_out[33] _1333__246/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_161_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1214__A _1247_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_22_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1816 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0992_ VGND VPWR _0993_/C _0992_/B _0992_/A _0992_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_18_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1475_ VGND VPWR _1475_/X _1475_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_141_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_613 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_545 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input91_A wbs_dat_i[27] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1110__C _1118_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_204_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_784 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output178_A _1483_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_174_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_799 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1119__A _1141_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_68_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_hold2_A hold2/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_123_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1260_ VGND VPWR _1255_/X _1254_/X _1256_/X _1260_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_211_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1191_ VGND VPWR _1188_/X _1187_/X _1189_/X _1191_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
Xinput8 VGND VPWR input8/X la_data_in[39] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_840 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0975_ _0975_/Y _0975_/B _0975_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_186_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0632__S _0636_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_31_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1458_ VGND VPWR _1458_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_19_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_615 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_790 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1339__252 irq[1] _1339__252/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_65_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0760_ _1118_/A _1478_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_200_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0691_ VPWR VGND _0986_/A _1491_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_155_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_780 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1312_ _1312_/Q _1241_/Y _1312_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_96_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1243_ VGND VPWR _1239_/X _1238_/X _1240_/X _1243_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_110_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1015__C _1065_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_211_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1174_ VGND VPWR _1171_/X _1169_/X _1173_/X _1174_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_65_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0958_ _0958_/B _0958_/X _1001_/A _0958_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_140_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0889_ _0889_/B _0889_/Y _0903_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_31_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput120 VPWR VGND io_oeb[19] _1456_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput131 VPWR VGND io_oeb[29] _1466_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput142 VPWR VGND io_oeb[5] _1442_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_118_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput153 VPWR VGND io_out[15] _1489_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_157_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput164 VPWR VGND io_out[25] _1499_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_138_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput175 VPWR VGND io_out[6] _1480_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput186 VPWR VGND la_data_out[16] _1490_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput197 VPWR VGND la_data_out[26] _1500_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_66_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1222__A _1246_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_102_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_327 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input54_A la_oenb[51] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_84_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0971__A _1141_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_91_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput11 VGND VPWR _1065_/B la_data_in[42] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0812_ _0812_/B _0822_/A _0812_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_204_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput22 VGND VPWR _0948_/C la_data_in[53] VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput33 VGND VPWR input33/X la_data_in[64] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput44 VGND VPWR _0814_/B la_oenb[41] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput55 VGND VPWR _0957_/A la_oenb[52] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0743_ VGND VPWR _1307_/D _0743_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput66 VGND VPWR _0819_/D la_oenb[63] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_171_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput77 input77/X wbs_dat_i[14] VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_116_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput88 VPWR VGND _0918_/C wbs_dat_i[24] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_192_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput99 VPWR VGND _1112_/A wbs_dat_i[5] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_196_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0674_ VGND VPWR _0674_/X _0674_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1226_ VGND VPWR _1223_/X _1222_/X _1224_/X _1226_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_6_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1157_ VPWR VGND hold2/X _1158_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1042__A _1486_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1310__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_164_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1088_ input8/X _1094_/C _1088_/A _1080_/A _1088_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__or4bb_4
XFILLER_0_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_687 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_514 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_410 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_658 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output160_A _1495_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_136_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1127__A _1127_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_45_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1011_ VGND VPWR _1031_/D _1025_/D _0938_/A _1013_/C _1489_/A _1070_/C VGND VPWR
+ sky130_fd_sc_hd__a41o_1
XFILLER_47_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0726_ VGND VPWR _0742_/S _1057_/B _1310_/Q _0727_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_172_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0657_ VGND VPWR _0665_/S _1323_/Q _0914_/A _0658_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_154_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0876__A _1080_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_58_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1209_ VGND VPWR _1204_/X _1203_/X _1205_/X _1209_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_66_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1500__A _1500_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0779__A1 _1132_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_166_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_834 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_551 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input17_A la_data_in[48] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_63_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_779 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_240 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_251 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_262 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_433 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1491_ VGND VPWR _1491_/X _1491_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_160 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_0_counter.clk_A _1152_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_94_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0630__A0 _1503_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_148_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0709_ VGND VPWR _0709_/X _0709_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1372__285 la_data_out[63] _1372__285/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input9_A la_data_in[40] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_98_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1230__A _1246_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_959 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_653 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1828 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0991_ _1491_/A _0992_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_14_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1356__269 la_data_out[47] _1356__269/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_86_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1474_ VGND VPWR _1474_/X _1474_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_140_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0873__B _1078_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_184_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1050__A _1050_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_36_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_636 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input84_A wbs_dat_i[20] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_128_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_796 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0958__B _0958_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_122_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1190_ VGND VPWR _1188_/X _1187_/X _1189_/X _1190_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_7_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput9 VGND VPWR input9/X la_data_in[40] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1086__B1 _1005_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0833__B1 _0832_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0974_ _0973_/X _0824_/X _0972_/Y _0990_/D input20/X _0975_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41oi_4
XFILLER_146_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1457_ VGND VPWR _1457_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1045__A _1111_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0884__A _0884_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_82_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_411 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_549 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1378__291 la_data_out[69] _1378__291/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_151_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0794__A _1502_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_150_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_811 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_71 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_82 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0690_ VGND VPWR _1317_/D _0690_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_170_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0969__A _0993_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_174_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1311_ _1311_/Q _1237_/Y _1311_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_135_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_792 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1242_ VGND VPWR _1239_/X _1238_/X _1240_/X _1242_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_38_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1173_ VPWR VGND _1205_/A _1173_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0957_ _0957_/A _0957_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_203_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0888_ _0888_/A _0903_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_173_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput110 VPWR VGND io_oeb[0] _1437_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_134_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput121 VPWR VGND io_oeb[1] _1438_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_192_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput132 VPWR VGND io_oeb[2] _1439_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_86_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput143 VPWR VGND io_oeb[6] _1443_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput154 VPWR VGND io_out[16] _1490_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput165 VPWR VGND io_out[26] _1500_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_153_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput176 VPWR VGND io_out[7] _1481_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_138_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput187 VPWR VGND la_data_out[17] _1491_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_142_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput198 VPWR VGND la_data_out[27] _1501_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_43_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1412__325 la_data_out[103] _1412__325/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_9_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1503__A _1503_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_83_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input47_A la_oenb[44] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1003 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1132__B _1132_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0811_ _0811_/C _0811_/B _0812_/B _0811_/D _0811_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_198_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput12 VGND VPWR _1055_/B la_data_in[43] VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput23 VGND VPWR _0941_/C la_data_in[54] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput34 la_data_in[65] hold2/A VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
Xinput45 VGND VPWR _0814_/C la_oenb[42] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0742_ VGND VPWR _0742_/S _1050_/A _1307_/Q _0743_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput56 VGND VPWR _0816_/B la_oenb[53] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_873 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xinput67 VGND VPWR _1151_/S la_oenb[64] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_155_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput78 wbs_dat_i[15] _1018_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_171_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput89 wbs_dat_i[25] _0907_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_116_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0673_ VGND VPWR _0692_/S _1320_/Q _0951_/A _0674_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_192_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1345 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1225_ VGND VPWR _1223_/X _1222_/X _1224_/X _1225_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_65_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1156_ _1473_/A _1156_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
XFILLER_65_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1087_ _1274_/D _1041_/X _1082_/Y _1062_/A _1086_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_41_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1489 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0881__B _0881_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_94_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_537 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_400 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input101_A wbs_dat_i[7] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_411 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_422 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1285__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output153_A _1489_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_105_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1143__A _1143_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_47_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1010_ VPWR VGND _1025_/D _1030_/A _1010_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_130_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0982__A _0982_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_408 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_482 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0725_ VGND VPWR _0725_/X _0725_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_155_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0656_ VPWR VGND _0914_/A _1498_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_171_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1153 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1208_ VGND VPWR _1204_/X _1203_/X _1205_/X _1208_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_150_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1139_ _1475_/A _1140_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_81_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1264 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_419 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1275 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_920 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1418__331 la_data_out[109] _1418__331/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_134_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_780 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_241 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_252 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_263 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_285 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_296 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1490_ VGND VPWR _1490_/X _1490_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1300__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_165_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0942__A2 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1 hold1/A hold1/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_39_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_807 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0708_ VGND VPWR _0717_/S _1313_/Q _1010_/A _0709_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_89_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0933__A2 input87/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_172_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0639_ VGND VPWR _0639_/S _1326_/Q _0891_/A _0640_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_67_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_260 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_counter.clk clkbuf_3_5_0_counter.clk/A _1296_/CLK VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_190_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0797__A _1481_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_46_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_687 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1140__B _1140_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_204_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0990_ _0990_/D _0990_/C _1142_/B _0990_/Y _0817_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_2
XFILLER_32_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1473_ VGND VPWR _1473_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_114_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0900__A2_N _0884_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_140_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1050__B _1050_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_580 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input77_A wbs_dat_i[14] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_136_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_495 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1086__A1 _1026_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_75_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0973_ _1001_/A _0973_/B _1092_/B _0973_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_146_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1456_ VGND VPWR _1456_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0884__B _0888_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_82_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1061__A _1125_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_517 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_823 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_856 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_72 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_83 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1310_ _1310_/Q _1236_/Y _1310_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_123_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0751__A0 _1102_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_173_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1241_ VGND VPWR _1239_/X _1238_/X _1240_/X _1241_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_77_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1172_ _1205_/A _1256_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_64_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0956_ _1287_/D _0869_/X _0954_/Y _0936_/Y _0955_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_146_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0887_ VGND VPWR _0831_/Y _0885_/Y _1067_/A _0887_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_31_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput111 VPWR VGND io_oeb[10] _1447_/X VGND VPWR sky130_fd_sc_hd__buf_2
XANTENNA__0879__B _0879_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xoutput122 VPWR VGND io_oeb[20] _1457_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput133 VPWR VGND io_oeb[30] _1467_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_192_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput144 VPWR VGND io_oeb[7] _1444_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_173_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput155 VPWR VGND io_out[17] _1491_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput166 VPWR VGND io_out[27] _1501_/A VGND VPWR sky130_fd_sc_hd__buf_2
XANTENNA__1056__A _1056_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xoutput177 VPWR VGND io_out[8] _1482_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_153_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput188 VPWR VGND la_data_out[18] _1492_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput199 VPWR VGND la_data_out[28] _1502_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_101_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1439_ VGND VPWR _1439_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_56_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1015 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_664 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0810_ _0810_/C _0810_/B _0812_/A _1088_/A _0810_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_204_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput13 VGND VPWR _1048_/C la_data_in[44] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput24 VGND VPWR _0932_/C la_data_in[55] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_7_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput35 VPWR VGND _0811_/A la_oenb[32] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_204_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput46 VGND VPWR _0814_/D la_oenb[43] VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1394__307 la_data_out[85] _1394__307/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_0741_ VGND VPWR _0741_/X _0741_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput57 VGND VPWR _0816_/C la_oenb[54] VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput68 VPWR VGND hold3/A la_oenb[65] VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_115_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_885 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xinput79 VPWR VGND _1001_/C wbs_dat_i[16] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_155_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0672_ _1047_/A _0692_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_170_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1435__348 la_data_out[126] _1435__348/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_83_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0724__A0 _1057_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1224_ VPWR VGND _1248_/A _1224_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1155_ _1156_/A _1256_/A _1255_/A hold2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_20_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_439 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1086_ _1026_/A _1005_/X _1086_/Y _1085_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0939_ _0940_/B _0962_/D _0936_/Y _0971_/D _0935_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31ai_1
XFILLER_147_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_549 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_412 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_423 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0954__B1 _0948_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_113_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0982__B _0982_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_494 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0724_ VGND VPWR _0744_/S _1310_/Q _1057_/B _0725_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_155_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0655_ VGND VPWR _1324_/D _0655_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_131_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1207_ VGND VPWR _1204_/X _1203_/X _1205_/X _1207_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_72_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1138_ _1268_/D _1027_/X _1136_/Y _1132_/A _1137_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__0892__B _0897_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_25_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1069_ _1483_/A _1070_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_41_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1298 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_814 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_910 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_220 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_264 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_286 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xhold2 hold2/X hold2/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_94_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0993__A _0997_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_54_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0707_ _1010_/A _1488_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_171_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0638_ _0891_/A _1501_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1275__CLK _1279_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1239__A _1247_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_5_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0797__B _1480_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_699 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input22_A la_data_in[53] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_36_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_265 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1298__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1022__C1 _1021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_5_961 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1472_ VGND VPWR _1472_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_140_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_941 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1034__D _1034_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1059__A _1067_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_526 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_386 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1002 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_821 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1649 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0990__B _1142_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_507 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0972_ _0972_/A _0972_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1362__275 la_data_out[53] _1362__275/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_105_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1455_ VGND VPWR _1455_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1313__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_209_771 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1061__B _1475_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_651 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1068__A2 _1065_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_27_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_835 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_868 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1346__259 la_data_out[37] _1346__259/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_73 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_84 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_562 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output176_A _1481_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_136_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1240_ VPWR VGND _1248_/A _1240_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1171_ VPWR VGND _1204_/A _1171_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0955_ _0929_/X _0910_/X _0955_/Y _0951_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_203_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0886_ VPWR VGND _1067_/A _1027_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_146_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput112 VPWR VGND io_oeb[11] _1448_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_86_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput123 VPWR VGND io_oeb[21] _1458_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput134 VPWR VGND io_oeb[31] _1468_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput145 VPWR VGND io_oeb[8] _1445_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_82_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput156 VPWR VGND io_out[18] _1492_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_192_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput167 VPWR VGND io_out[28] _1502_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput178 VPWR VGND io_out[9] _1483_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_153_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput189 VPWR VGND la_data_out[19] _1493_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0742__A1 _1050_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_25_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1438_ VGND VPWR _1438_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1072__A _1072_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_210_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_243 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_265 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_809 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1247__A _1247_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_536 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1027 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput14 VGND VPWR _1034_/C la_data_in[45] VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput25 VPWR VGND la_data_in[56] _0920_/C VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0740_ VGND VPWR _0744_/S _1307_/Q _1050_/A _0741_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput36 VGND VPWR _0811_/B la_oenb[33] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput47 VGND VPWR _0813_/A la_oenb[44] VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput58 VGND VPWR _0816_/D la_oenb[55] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_183_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput69 VPWR VGND _0787_/A la_oenb[66] VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_170_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0671_ VPWR VGND _1047_/A _0897_/B VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_100_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1157__A hold2/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_170_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1223_ VPWR VGND _1247_/A _1223_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1336 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1369 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1154_ hold3/X input70/X _1256_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2b_4
XFILLER_20_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1085_ _1115_/D _1125_/A _1085_/X _1132_/A _1085_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_94_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1368__281 la_data_out[59] _1368__281/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1107__A1_N _0832_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_178_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0938_ _0938_/A _0971_/D _0992_/B _0961_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_2
XFILLER_159_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0869_ _0869_/X _1097_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0715__A1 _1030_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_402 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_690 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_801 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0954__A1 _0944_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_138_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input52_A la_oenb[49] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_65_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1440__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_62_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1402__315 la_data_out[93] _1402__315/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_198_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0723_ _1047_/A _0744_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_155_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0654_ VGND VPWR _0663_/S _0888_/A _1324_/Q _0655_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_170_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1206_ VGND VPWR _1204_/X _1203_/X _1205_/X _1206_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_6_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1137_ _1100_/Y _0861_/X _1137_/Y _1115_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_81_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1233 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1068_ _1066_/Y _1067_/Y _1276_/D _1064_/Y _1065_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_2
XFILLER_55_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1095 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1019 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_922 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_232 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_254 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_265 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1154__B hold3/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_94_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xhold3 VPWR VGND hold3/X hold3/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_94_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1170__A _1255_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0706_ VGND VPWR _1314_/D _0706_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_132_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0637_ VGND VPWR _1327_/D _0637_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1080__A _1080_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_65_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_903 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0797__C _1479_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_27_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1255__A _1255_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_66_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_678 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input15_A la_data_in[46] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_29_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_233 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1022__B1 _0861_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_114_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1471_ VGND VPWR _1471_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_114_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1408__321 la_data_out[99] _1408__321/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_63_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_538 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1059__B _1059_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_178_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input7_A la_data_in[38] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_376 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_475 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1135__D _1142_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0971_ _0971_/C _1000_/B _0975_/A _0971_/D _1141_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_38_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0999__A _1050_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_69_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_counter.clk clkbuf_0_counter.clk/X _1152_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_58_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_781 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1454_ VGND VPWR _1454_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_663 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1288__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_302 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1385__298 la_data_out[76] _1385__298/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XPHY_52 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_74 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_96 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_981 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input82_A wbs_dat_i[19] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_128_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output169_A _1476_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_155_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1443__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_113_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1170_ _1204_/A _1255_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_37_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0954_ _0944_/Y _1000_/B _0954_/Y _0953_/Y _0948_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_1
XFILLER_146_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0885_ _0885_/B _0885_/Y _0889_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_88_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput113 VPWR VGND io_oeb[12] _1449_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_12_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput124 VPWR VGND io_oeb[22] _1459_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_115_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput135 VPWR VGND io_oeb[32] _1469_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_177_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput146 VPWR VGND io_oeb[9] _1446_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput157 VPWR VGND io_out[19] _1493_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_82_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput168 VPWR VGND io_out[29] _1503_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_192_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput179 VPWR VGND la_data_out[0] _1474_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_86_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1437_ VGND VPWR _1437_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1299_ _1299_/Q _1219_/Y _1299_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_56_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_165 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_198 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput15 VGND VPWR _1021_/C la_data_in[46] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_167_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput26 VPWR VGND la_data_in[57] input26/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput37 VGND VPWR _0811_/C la_oenb[34] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1438__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_128_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput48 VGND VPWR _0813_/B la_oenb[45] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_865 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xinput59 VPWR VGND la_oenb[56] _0820_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1303__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_0670_ VPWR VGND _0951_/A _1495_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_183_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1173__A _1205_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_65_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1222_ VPWR VGND _1246_/A _1222_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1153_ _1255_/A hold3/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_93_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1084_ _1115_/D _1132_/C _1132_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_20_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1222 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0937_ _0950_/A _0962_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_159_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0868_ _1027_/A _1097_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__1067__B _1067_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_162_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0799_ _0901_/A _0985_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_153_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1083__A _1125_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_88_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_909 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_403 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_414 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_625 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_485 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_389 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input45_A la_oenb[42] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_171_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1168__A hold2/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_129_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0722_ _1057_/B _1485_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_200_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0653_ VGND VPWR _0653_/X _0653_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0800__A _1486_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1145 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1205_ VPWR VGND _1205_/A _1205_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_211_1189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_205 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1136_ _1136_/Y _1136_/A _1136_/C _1136_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_65_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1067_ _1067_/B _1067_/Y _1067_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_41_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1289 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_827 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1009 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1425__338 la_data_out[116] _1425__338/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_73_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_934 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_244 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_255 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0624__A1 _1505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_73_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_266 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_288 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output151_A _1487_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1451__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_208_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0705_ VGND VPWR _0715_/S _1489_/A _1314_/Q _0706_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_171_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0636_ VGND VPWR _0636_/S _1502_/A _1327_/Q _0637_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_63_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1119_ _1122_/A _1141_/A _1119_/C _1141_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_26_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_915 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0797__D _1478_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_27_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1098__A1 _1088_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_28_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1022__A1 _1016_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_153_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1446__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_99_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1470_ VGND VPWR _1470_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_153_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1181__A _1205_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_209_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0836__A1 _0841_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_63_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0836__B2 _0877_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_208_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_629 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0619_ _1021_/B _0639_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_594 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_204 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_955 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_487 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_333 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0970_ _0970_/B _0971_/C _0970_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_105_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1453_ VGND VPWR _1453_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1081 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_336 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_64 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_86 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_97 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input75_A wbs_dat_i[12] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1608 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0953_ _0953_/Y _0953_/A _0997_/A _0993_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_202_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0803__A _1493_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_70_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0884_ _0885_/B _0888_/A _0884_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_185_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput114 VPWR VGND io_oeb[13] _1450_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput125 VPWR VGND io_oeb[23] _1460_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_115_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput136 VPWR VGND io_oeb[33] _1470_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput147 VPWR VGND io_out[0] _1474_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_173_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput158 VPWR VGND io_out[1] _1475_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1505_ VGND VPWR _1505_/X _1505_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xoutput169 VPWR VGND io_out[2] _1476_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_115_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1298_ _1298_/Q _1218_/Y _1298_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_110_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_601 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_634 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1352__265 la_data_out[43] _1352__265/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_59_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_counter.clk clkbuf_0_counter.clk/X clkbuf_2_1_0_counter.clk/A VGND VPWR
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_169_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_100 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_634 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_790 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput16 VPWR VGND la_data_in[47] _1015_/B VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput27 VGND VPWR _0897_/C la_data_in[58] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_167_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput38 VGND VPWR _0811_/D la_oenb[35] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_183_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput49 VGND VPWR _0813_/C la_oenb[46] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_182_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1454__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_174_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1221_ VGND VPWR _1214_/X _1212_/X _1216_/X _1221_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_84_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1152_ VGND VPWR _1152_/X _1152_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_37_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1083_ _1125_/B _1132_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_53_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1289 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0936_ _0951_/A _0936_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_88_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0867_ _0862_/Y _0866_/Y _1295_/D _0795_/B _0790_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22ai_1
XFILLER_146_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0798_ _1062_/D _0901_/A _1077_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_192_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1278__CLK _1279_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_130_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1336__249 io_out[36] _1336__249/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_170_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1872 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_404 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_415 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input38_A la_oenb[35] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_66_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1116__B1 _1005_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_59_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0618__A _0897_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1449__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_106_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0721_ VGND VPWR _1311_/D _0721_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_129_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0652_ VGND VPWR _0665_/S _1324_/Q _0888_/A _0653_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_170_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0800__B _1485_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_170_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1204_ VPWR VGND _1204_/A _1204_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1168 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1135_ _1142_/D input3/X _1135_/B _1136_/C _0811_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_93_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1066_ input73/X _0790_/A _1066_/Y _1079_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_20_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0919_ _1073_/B _1080_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_162_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1094__A _1094_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_153_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_212 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_234 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_946 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_256 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_267 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1358__271 la_data_out[49] _1358__271/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_101_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0993__D _0993_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_208_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_counter.clk clkbuf_3_1_0_counter.clk/A _1316_/CLK VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__1179__A _1203_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_34_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0704_ VGND VPWR _0704_/X _0704_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0811__A _0811_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_144_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0635_ VGND VPWR _0635_/X _0635_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_131_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1316__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_39_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1118_ _1118_/B _1119_/C _1118_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_81_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1049_ _1049_/Y _1049_/A _1049_/C _1049_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_41_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1089__A _1477_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_70_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_703 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1022__A2 input77/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_201_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_953 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0777__S _1034_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_151_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1462__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_136_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_680 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_933 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_977 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0836__A2 _0945_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_63_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0772__A1 _1125_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_132_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0618_ _1021_/B _0897_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_63_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1149 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0763__A1 _1118_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_146_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_967 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_207 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input20_A la_data_in[51] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_188_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_389 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1457__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_199_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1452_ VGND VPWR _1452_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_65 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_87 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_98 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_569 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input68_A la_oenb[65] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_151_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0736__A1 _1059_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_194_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0883__A1_N _0869_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_53_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0952_ _0997_/A _0952_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_32_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0883_ _1294_/D _0869_/X _0881_/Y _0882_/Y _0873_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__0803__B _1492_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_88_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1187__A _1203_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_200_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput115 VPWR VGND io_oeb[14] _1451_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput126 VPWR VGND io_oeb[24] _1461_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput137 VPWR VGND io_oeb[34] _1471_/X VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput148 VPWR VGND io_out[10] _1484_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1504_ VGND VPWR _1504_/X _1504_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xoutput159 VPWR VGND io_out[20] _1494_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1297_ _1505_/A _1217_/Y _1297_/D _1326_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_3_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_646 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput17 VGND VPWR _1002_/C la_data_in[48] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput28 VGND VPWR _0892_/C la_data_in[59] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xinput39 VGND VPWR _0810_/A la_oenb[36] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_377 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output174_A _1479_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_136_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1220_ VGND VPWR _1214_/X _1212_/X _1216_/X _1220_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_113_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1151_ VGND VPWR wb_clk_i input33/X _1151_/S _1152_/A VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_93_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1470__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_168_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0893__B1 _0892_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_93_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1082_ _1082_/Y _1082_/A _1082_/C _1082_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_0_1406 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0935_ _1496_/A _0935_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_124_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0866_ VGND VPWR _0866_/Y _0865_/X _0873_/A _0849_/A _0863_/Y VGND VPWR sky130_fd_sc_hd__a31oi_1
XFILLER_106_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0797_ _1480_/A _1481_/A _1062_/D _1478_/A _1479_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4_2
XFILLER_115_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1375__288 la_data_out[66] _1375__288/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_130_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_405 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_837 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1116__A1 _1100_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0720_ VGND VPWR _0742_/S _1486_/A _1311_/Q _0721_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_200_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0651_ _0888_/A _1499_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_7_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1465__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_143_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0800__C _1484_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_174_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1203_ VPWR VGND _1203_/A _1203_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1134_ _1136_/B _1134_/B _1134_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_53_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_793 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1065_ _0814_/C _1065_/Y _1065_/B _1065_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3b_4
XFILLER_209_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_457 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1078__C _1078_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_159_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0918_ _0918_/B _1094_/A _0921_/B _1094_/C _0918_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4_2
XFILLER_198_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0849_ _0849_/A _0849_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_162_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1094__B _1094_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_68_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_719 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_213 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_224 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_257 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input50_A la_oenb[47] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_152_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_177 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1268__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_206_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0703_ VGND VPWR _0717_/S _1314_/Q _1489_/A _0704_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_472 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1195__A _1203_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_144_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0634_ VGND VPWR _0639_/S _1327_/Q _1502_/A _0635_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_131_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1117_ _1271_/D _1041_/X _1114_/Y _1110_/B _1116_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_54_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1048_ _1121_/D _1048_/C _1073_/B _1049_/C _0813_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_110_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1089__B _1476_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_142_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1390__303 la_data_out[81] _1390__303/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_153_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1431__344 la_data_out[122] _1431__344/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_153_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_243 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input98_A wbs_dat_i[4] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_160_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_932 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_692 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0617_ _0897_/B _0854_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_131_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1415__328 la_data_out[106] _1415__328/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_63_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_445 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_803 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input13_A la_data_in[44] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_206_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1306__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_195_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1451_ VGND VPWR _1451_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_99_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1473__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_84_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_806 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input5_A la_data_in[36] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_86_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_66 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1329__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_99 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_962 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_526 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_809 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0951_ _0951_/B _0953_/A _0951_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_202_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1468__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0882_ _0849_/X _0848_/X _0882_/Y _0809_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XANTENNA__0803__C _1491_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_179_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput116 VPWR VGND io_oeb[15] _1452_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_56_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput127 VPWR VGND io_oeb[25] _1462_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput138 VPWR VGND io_oeb[35] _1472_/X VGND VPWR sky130_fd_sc_hd__buf_2
X_1503_ VGND VPWR _1503_/X _1503_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xoutput149 VPWR VGND io_out[11] _1485_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1296_ _1504_/A _1210_/Y _1296_/D _1296_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_209_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0663__A1 _1497_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1097__B _1481_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_197_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0654__A1 _0888_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_781 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1064__D1 _1078_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_54_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_864 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput18 VGND VPWR _0990_/C la_data_in[49] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_input80_A wbs_dat_i[17] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xinput29 VPWR VGND la_data_in[60] input29/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output167_A _1502_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_151_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1150_ _1146_/Y _1266_/D _1149_/X _1140_/B _1027_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1081_ _1121_/D input9/X _1135_/B _1082_/C _0814_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_19_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1418 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0934_ _0832_/X _1289_/D VGND VPWR _0933_/Y _0930_/Y _1497_/A VGND VPWR sky130_fd_sc_hd__a2bb2oi_1
XFILLER_72_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0865_ input93/X _0864_/X _0907_/A _0842_/X _0865_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_88_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0796_ _1477_/A _1474_/A _1475_/A _1476_/A _1077_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_200_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1279_ _1487_/A _1184_/Y _1279_/D _1279_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_71_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_406 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0636__A1 _1502_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_783 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0650_ VGND VPWR _1325_/D _0650_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0800__D _1483_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_98_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1481__A _1481_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_113_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1202_ VGND VPWR _1196_/X _1195_/X _1197_/X _1202_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_61_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1133_ _1136_/A _1141_/A _1133_/C _1141_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_26_709 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1064_ _1059_/Y _1062_/X _1078_/B _1063_/X _1078_/C _1064_/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_39_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1033 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0825__A _0834_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_209_1044 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1342__255 la_data_out[33] _1342__255/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_33_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0917_ _1094_/C _0917_/A _0917_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_159_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0848_ VPWR VGND _0848_/X _1005_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_161_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0779_ VGND VPWR _0785_/S _1132_/B _1300_/Q _0780_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__1094__C _1094_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0857__A1 _0848_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__0828__C_N _1094_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_79_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1793 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_797 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_247 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input43_A la_oenb[40] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_171_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_580 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_753 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0645__A _1500_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_952 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1476__A _1476_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_195_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0702_ VGND VPWR _1315_/D _0702_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_144_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0633_ VGND VPWR _1328_/D _0633_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_98_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1116_ _1100_/Y _1005_/X _1116_/Y _1115_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_148_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1047_ VPWR VGND _1121_/D _1047_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_734 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1089__C _1475_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_266 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_944 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0616_ _0854_/A _0834_/B _0834_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_193_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_358 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1348__261 la_data_out[39] _1348__261/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_41_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_914 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_925 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_848 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0907__B _0907_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_206_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1450_ VGND VPWR _1450_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_206_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_490 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_870 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1184 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1155__B1 _1256_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_86_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_67 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_974 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_996 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1146__B1 _0790_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_89_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0918__A _1094_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_65_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0950_ _0999_/B _0992_/A _0951_/B _0961_/C _0950_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_13_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0881_ _0881_/Y _0881_/B _0881_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_158_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0803__D _1490_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1484__A _1484_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_66_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput117 VPWR VGND io_oeb[16] _1453_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_127_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput128 VPWR VGND io_oeb[26] _1463_/X VGND VPWR sky130_fd_sc_hd__buf_2
X_1502_ VGND VPWR _1502_/X _1502_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xoutput139 VPWR VGND io_oeb[36] _1473_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1137__B1 _0861_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_68_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1295_ _1503_/A _1209_/Y _1295_/D _1296_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_3_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_counter.clk clkbuf_2_3_0_counter.clk/A clkbuf_3_7_0_counter.clk/A VGND
+ VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_865 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0738__A _1482_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_115_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input108_A wbs_stb_i VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_814 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_876 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput19 VGND VPWR input19/X la_data_in[50] VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input73_A wbs_dat_i[10] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_124_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1080_ VPWR VGND _1135_/B _1080_/A VGND VPWR sky130_fd_sc_hd__buf_4
XANTENNA__0893__A2 input91/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_168_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1479__A _1479_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_106 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0933_ _0933_/Y _0790_/A _1001_/A _0872_/B _0932_/X input87/X VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a311oi_4
XFILLER_174_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0864_ VGND VPWR _0897_/B _0864_/X _0819_/B _0864_/C VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_179_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0795_ _0795_/A _0809_/A _0795_/B _0873_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_114_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1319__CLK _1330_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1021 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1278_ _1486_/A _1183_/Y _1278_/D _1279_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_186_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1054 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_407 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1150__A1_N _1146_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_902 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_counter.clk_A clkbuf_0_counter.clk/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__0931__A _0982_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1201_ VGND VPWR _1196_/X _1195_/X _1197_/X _1201_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_66_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1132_ VGND VPWR _1133_/C _1132_/B _1132_/A _1132_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_4_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1063_ _1070_/C _1067_/B _1059_/B _1070_/A _1063_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_4_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1056 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1381__294 la_data_out[72] _1381__294/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_198_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0841__A _0841_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_0916_ _0830_/Y _0828_/X _0921_/A _0980_/A _0915_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_1
XFILLER_30_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0847_ _1005_/A _0861_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_198_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0778_ VGND VPWR _0778_/X _0778_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_115_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_204 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_242 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_226 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_237 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_248 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_647 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input36_A la_oenb[33] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0926__A _1493_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_798 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1365__278 la_data_out[56] _1365__278/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_206_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_964 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0701_ VGND VPWR _0715_/S _0993_/D _1315_/Q _0702_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_183_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0632_ VGND VPWR _0636_/S _1503_/A _1328_/Q _0633_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1492__A _1492_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_80_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1115_ _1132_/A _1115_/A _1115_/X _1125_/A _1115_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_93_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_529 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1046_ _1049_/B _1072_/B _1046_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_181_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_713 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_746 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1089__D _1474_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_52_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_80 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_606 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_978 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0656__A _1498_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_91_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1487__A _1487_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_34_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1029_ _1054_/C _1078_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_41_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_727 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0905__D1 _0980_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_131_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_241 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_970 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_981 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_882 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1421__334 la_data_out[112] _1421__334/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_34_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1010__A _1010_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_136_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1155__A1 hold2/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_68 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_953 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1091__B1 _1481_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_50_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1146__A1 _0980_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_624 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0657__A0 _0914_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_146_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1405__318 la_data_out[96] _1405__318/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_60_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0880_ _0879_/X _1142_/B _0874_/Y _0990_/D input29/X _0881_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41oi_4
XFILLER_201_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput118 VPWR VGND io_oeb[17] _1454_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_142_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput129 VPWR VGND io_oeb[27] _1464_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_182_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1501_ VGND VPWR _1501_/X _1501_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1137__A1 _1100_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_190_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1294_ _1502_/A _1208_/Y _1294_/D _1294_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_83_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0639__A0 _0891_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_210_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_321 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_826 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_888 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input66_A la_oenb[63] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_184_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0932_ VGND VPWR _0947_/A _0932_/X _0816_/D _0932_/C VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_163_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0863_ _0873_/D _0863_/Y _1503_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_179_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1495__A _1495_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_174_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0794_ _1502_/A _0873_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_127_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1277_ _1485_/A _1182_/Y _1277_/D _1281_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_84_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1427__340 la_data_out[118] _1427__340/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XPHY_419 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_468 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0749__A _1480_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_82_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_914 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output172_A _1477_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_67_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1200_ VGND VPWR _1196_/X _1195_/X _1197_/X _1200_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_61_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1131_ _1269_/D _1027_/X _1129_/Y _1125_/A _1130_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_187_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1062_ _1062_/C _1062_/A _1062_/X _1125_/A _1062_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_0_1217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1239 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1028__B1 _1010_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0915_ _0915_/X _0922_/B _0992_/A _0992_/B _0915_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_120_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0846_ _0833_/Y _0790_/X _0845_/Y _1505_/A _1297_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_4
XFILLER_175_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0777_ VGND VPWR _1034_/D _1300_/Q _1132_/B _0778_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1329_ _1329_/Q _1264_/Y _1329_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_25_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1740 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1751 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_205 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_238 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_659 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input29_A la_data_in[60] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_207_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0926__B _0979_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_74_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_766 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1309__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_160_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_420 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0700_ VGND VPWR _0700_/X _0700_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_976 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_464 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0631_ VGND VPWR _0631_/X _0631_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1114_ _1114_/Y _1114_/A _1114_/C _1114_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_4_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1045_ _1049_/A _1111_/A _1045_/C _1078_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_53_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1013__A _1078_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_39_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0829_ _0841_/A _0907_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_780 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1332__245 io_out[32] _1332__245/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_125_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0937__A _0950_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_23_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0956__A1_N _0869_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_189_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0672__A _1047_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_784 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_261 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1028_ _1022_/Y _1280_/D _1026_/Y _1027_/X _1010_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_210_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_828 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0684__A1 _1493_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_79_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input96_A wbs_dat_i[31] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_264 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0675__A1 _0951_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_75_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1498__A _1498_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_182_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1010__B _1030_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_125_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1155__A2 _1255_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_99_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_910 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1091__A1 _1102_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_23_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_396 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0918__C _0918_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_66_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_636 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_102 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input11_A la_data_in[42] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_79_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1111__A _1111_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_207_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0950__A _0950_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_16_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_367 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_540 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1500_ VGND VPWR _1500_/X _1500_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xoutput119 VPWR VGND io_oeb[18] _1455_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_126_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1338__251 irq[0] _1338__251/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_99_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1293_ _1501_/A _1207_/Y _1293_/D _1296_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_81_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0860__A _1502_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_34_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input3_A la_data_in[34] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_86_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0920__D _1034_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_108_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input59_A la_oenb[56] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_97_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0945__A _0982_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0931_ _1001_/A _0982_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_92_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0862_ _0849_/X _0861_/X _0862_/Y _0860_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_35_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0793_ _1503_/A _0795_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_157_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1016__A _1094_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1276_ _1484_/A _1178_/Y _1276_/D _1281_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_186_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_361 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1877 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1888 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_753 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_439 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_613 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output165_A _1500_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_863 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1107 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1130_ _1100_/Y _0861_/X _1130_/Y _1062_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_66_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1061_ _1062_/C _1125_/B _1132_/C _1475_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_4_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1028__B2 _1027_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_159_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0914_ _0914_/A _0915_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_72_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0845_ _0840_/X _0844_/X _0845_/Y _0849_/A _0873_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_2
XFILLER_88_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0776_ VPWR VGND _1034_/D _0877_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_200_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1328_ _1328_/Q _1263_/Y _1328_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_29_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1259_ VGND VPWR _1255_/X _1254_/X _1256_/X _1259_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_77_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_756 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_239 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_277 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0926__C _1491_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_16_712 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_778 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0630_ VGND VPWR _0639_/S _1328_/Q _1503_/A _0631_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_109_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1113_ _1121_/D input6/X _1135_/B _1114_/C _0810_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_187_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1044_ _1045_/C _1070_/C _1070_/A _1044_/B _1050_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_39_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1013__B _1013_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_39_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0828_ _0917_/A _0917_/B _1094_/A _0828_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
XFILLER_89_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0759_ VGND VPWR _1304_/D _0759_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1204__A _1204_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_38_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1560 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_748 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input41_A la_oenb[38] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_641 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1371__284 la_data_out[62] _1371__284/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_88_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_949 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1100__B1 _1080_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_796 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0863__A _1503_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1027_ VPWR VGND _1027_/X _1027_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_53_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1355__268 la_data_out[46] _1355__268/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_115_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input89_A wbs_dat_i[25] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_200_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1149__B1 _1148_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1109__A _1109_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_181_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0918__D _1094_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1271__CLK _1279_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_44_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_counter.clk clkbuf_3_7_0_counter.clk/A _1279_/CLK VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_198_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1377__290 la_data_out[68] _1377__290/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_9_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1292_ _1500_/A _1206_/Y _1292_/D _1296_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_42_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1021__B _1021_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_31_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0860__B _0922_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_140_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1040__A1_N _0966_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1294__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_114_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_423 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1212__A _1246_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_208_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_802 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1088__C_N _1080_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_96_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1411__324 la_data_out[102] _1411__324/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_133_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_401 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0945__B _0945_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_189_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0961__A _1070_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_0930_ _1497_/A _0927_/X _0930_/Y _0929_/X _0922_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_1
XFILLER_42_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0861_ VPWR VGND _0861_/X _0861_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_158_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0792_ _1504_/A _0795_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_31_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1016__B _1016_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_28_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1275_ _1483_/A _1177_/Y _1275_/D _1279_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_68_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0855__B _0947_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_37_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1032__A _1111_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_52_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_632 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_308 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input106_A wbs_sel_i[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_151_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0781__A _1474_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_208_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_643 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input71_A wbs_cyc_i VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_171_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output158_A _1475_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_191_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0720__A1 _1486_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1060_ _1477_/A _1125_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_207_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1004 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_908 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_407 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0691__A _1491_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1002__D _1034_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_174_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0913_ _0985_/A _0992_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_119_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0844_ input96/X _0843_/X _0918_/B _0842_/X _0844_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_11_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0775_ VPWR VGND _0877_/A _0854_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_66_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1327_ _1327_/Q _1262_/Y _1327_/D _1330_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_211_1631 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1653 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1258_ VGND VPWR _1255_/X _1254_/X _1256_/X _1258_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_186_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1189_ VPWR VGND _1205_/A _1189_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1775 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0776__A _0877_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_130_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0926__D _1490_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_210_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_650 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1417__330 la_data_out[108] _1417__330/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_180_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_160 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0686__A _1492_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_120_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1112_ _1114_/B _1143_/B _1112_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_43_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_551 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1043_ VGND VPWR _1050_/C _1484_/A _1057_/B _1483_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_4_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0827_ VPWR VGND _1094_/A _0834_/C VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_176_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0758_ VGND VPWR _0767_/S _1109_/A _1304_/Q _0759_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_143_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0689_ VGND VPWR _0689_/S _0979_/A _1317_/Q _0690_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1461 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1572 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0620__A0 _1505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_138_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input34_A la_data_in[65] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0687__A0 _0979_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_521 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1100__A1 _1094_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1100__B2 _0947_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_43_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0678__A0 _0950_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1026_ _1026_/Y _1026_/A _1026_/C _1026_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_39_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1215__A _1256_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_69_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_557 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_517 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1149__B2 _0811_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_141_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0948__B _1142_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_114_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_995 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1019__B _1489_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_144_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1009_ _1031_/D _1484_/A _1486_/A _1485_/A _1483_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_23_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_888 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_989 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_538 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_counter.clk clkbuf_2_1_0_counter.clk/A clkbuf_3_1_0_counter.clk/A VGND
+ VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_173_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1291_ _1499_/A _1202_/Y _1291_/D _1296_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_81_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1489_ VGND VPWR _1489_/X _1489_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_619 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1250 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0860_ _0922_/B _0922_/A _0860_/Y _0860_/D _1502_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_35_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0791_ _1298_/Q _0790_/X _0636_/S _1298_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_10_891 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1016__C _1094_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1274_ _1482_/A _1176_/Y _1274_/D _1279_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_42_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0628__S _0636_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_83_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0989_ _0989_/A _0989_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_69_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1393__306 la_data_out[84] _1393__306/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_175_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1434__347 la_data_out[125] _1434__347/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_114_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1223__A _1247_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_76_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input64_A la_oenb[61] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1133__A _1141_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_130_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_419 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1284__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_187_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0912_ _1291_/D _0869_/X _0909_/Y _0903_/D _0911_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_50_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0843_ _0819_/D _0843_/X _0843_/C _0877_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_50_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0774_ _1475_/A _1132_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_157_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1326_ _1326_/Q _1261_/Y _1326_/D _1326_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_9_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1643 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1007__A1_N _0966_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1257_ VGND VPWR _1255_/X _1254_/X _1256_/X hold1/A VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_84_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1043__A _1057_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_37_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1188_ VPWR VGND _1204_/A _1188_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1765 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_208 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1787 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_452 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0831__A1_N _1021_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_49_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_736 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0792__A _1504_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_55_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_706 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output170_A _1504_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_197_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0967__A _0997_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_79_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1111_ _1114_/A _1111_/A _1111_/C _1141_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_43_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1042_ _1486_/A _1044_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_207_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0826_ _0834_/B _0917_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_190_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0757_ VGND VPWR _0757_/X _0757_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0688_ VGND VPWR _0688_/X _0688_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0877__A _0877_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_170_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1309_ _1309_/Q _1235_/Y _1309_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1501__A _1501_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_1584 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1399__312 la_data_out[90] _1399__312/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_40_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_621 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0787__A _0787_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_125_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input27_A la_data_in[58] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_87_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1114__C _1114_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0953__C _0997_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_204_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1322__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_176_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_297 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0697__A _1490_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_98_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1025_ _1031_/D _1050_/B _1026_/C _1025_/D _1050_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XANTENNA__0636__S _0636_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_35_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0809_ _0809_/B _0809_/Y _0809_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_85_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_429 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1231__A _1247_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_57_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1125__B _1125_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_759 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_853 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1141__A _1141_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_127_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0980__A _0980_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_207_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_380 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1089 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1008_ _1077_/A _1070_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_300 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0890__A _1500_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_91_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1361__274 la_data_out[52] _1361__274/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_41_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_237 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input94_A wbs_dat_i[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_554 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1290_ _1498_/A _1201_/Y _1290_/D _1296_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_209_501 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_209 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1345__258 la_data_out[36] _1345__258/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_189_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1046__A _1046_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_59_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1488_ VGND VPWR _1488_/X _1488_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_815 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_798 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_347 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1122__C _1122_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_37_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0790_ VPWR VGND _0790_/X _0790_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_881 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1273_ _1481_/A _1175_/Y _1273_/D _1281_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_81_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1836 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_678 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0988_ _1284_/D _0966_/X _0984_/Y _0980_/D _0987_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_140_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input1_A la_data_in[32] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_86_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1504__A _1504_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_68_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_745 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1367__280 la_data_out[58] _1367__280/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_19_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_573 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input57_A la_oenb[54] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_78_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_244 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1130__B1 _0861_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_59_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0911_ _0849_/X _0910_/X _0911_/Y _0889_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_147_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0842_ VPWR VGND _0945_/B _0842_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0773_ VGND VPWR _1301_/D _0773_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1325_ _1325_/Q _1260_/Y _1325_/D _1326_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_29_509 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1256_ VGND VPWR _1256_/X _1256_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_83_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1666 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1043__B _1484_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_168_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1187_ VPWR VGND _1203_/A _1187_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_409 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1799 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1401__314 la_data_out[92] _1401__314/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_608 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_258 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_718 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_925 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output163_A _1498_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_158_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1110_ VGND VPWR _1111_/C _1110_/B _1110_/A _1118_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_43_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1041_ _1097_/A _1041_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_24_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1103__B1 _1480_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_34_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_781 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0825_ _0834_/A _0917_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_176_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0756_ VGND VPWR _0770_/S _1304_/Q _1109_/A _0757_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_66_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0687_ VGND VPWR _0692_/S _1317_/Q _0979_/A _0688_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_66_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1054__A _1078_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_22_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1308_ _1308_/Q _1234_/Y _1308_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_211_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1239_ VPWR VGND _1247_/A _1239_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0908__B1 _0907_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_49_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_633 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1274__CLK _1279_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_94_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1139__A _1475_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_171_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0978__A _0986_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_28_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1024_ VGND VPWR _1050_/B _1031_/D _1050_/A _1026_/B _1010_/A _1030_/A VGND VPWR
+ sky130_fd_sc_hd__a41o_1
XFILLER_39_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0808_ _0949_/A _0985_/A _0809_/B _0860_/D _0922_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4_2
XFILLER_146_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0888__A _0888_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_143_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0739_ VPWR VGND _1050_/A _1077_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_46_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_854 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1407__320 la_data_out[98] _1407__320/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_25_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1382 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_430 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0948__D _1142_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1125__C _1132_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_392 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1035__C _1035_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_210_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1057 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1007_ _1282_/D _0966_/X _1003_/Y _0999_/C _1006_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_35_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1312__CLK _1316_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_122_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_824 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input87_A wbs_dat_i[23] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_750 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1152__A _1152_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_188_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0991__A _1491_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__1058__A2 _1055_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_51_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1384__297 la_data_out[75] _1384__297/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_149_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1487_ VGND VPWR _1487_/X _1487_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_113_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_827 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_921 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_965 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0986__A _0986_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_150_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1272_ _1480_/A _1174_/Y _1272_/D _1281_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_133_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1733 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_657 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0987_ _0929_/X _0910_/X _0987_/Y _0986_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_101_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_552 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0705__A1 _1489_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_78_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1130__A1 _1100_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_37_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0910_ _1005_/A _0910_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_53_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0841_ _0841_/A _0918_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0772_ VGND VPWR _0785_/S _1125_/B _1301_/Q _0773_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1324_ _1324_/Q _1259_/Y _1324_/D _1326_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_111_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1255_ VPWR VGND _1255_/A _1255_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_204_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1043__C _1483_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_42_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1186_ VGND VPWR _1180_/X _1179_/X _1181_/X _1186_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_209_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0880__B1 _0879_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_16_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_865 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput240 VPWR VGND wbs_dat_o[6] _0752_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_160_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_581 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0699__A0 _0993_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_47_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input104_A wbs_sel_i[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_71_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output156_A _1492_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_78_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1144__B _1144_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_130_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1040_ _1279_/D _0966_/X _1035_/Y _1031_/B _1039_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_130_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0862__B1 _0861_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_146_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1424__337 la_data_out[115] _1424__337/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_148_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0824_ VPWR VGND _0824_/X _0824_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_11_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_813 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_970 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0755_ _1109_/A _1479_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_102_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0686_ VPWR VGND _0979_/A _1492_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_118_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1307_ _1307_/Q _1233_/Y _1307_/D _1316_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_29_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1453 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1238_ VPWR VGND _1246_/A _1238_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1070__A _1070_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1169_ VPWR VGND _1203_/A _1169_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1597 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_417 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_656 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_513 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0844__B1 _0843_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_108_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0978__B _1490_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_124_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1023_ _0958_/C _1021_/B _1016_/B _0824_/X _1026_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a22oi_4
XFILLER_35_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0807_ _0860_/D _1499_/A _1501_/A _1500_/A _1498_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_50_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0738_ VPWR VGND _1482_/A _1077_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0669_ VGND VPWR _1321_/D _0669_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_39_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_893 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1394 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_549 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_665 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_910 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_442 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input32_A la_data_in[63] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1114 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_433 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_360 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_371 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_382 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1389__302 la_data_out[80] _1389__302/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
Xclkbuf_3_3_0_counter.clk clkbuf_3_3_0_counter.clk/A _1330_/CLK VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_66_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1069 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_192 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1006_ _0929_/X _1005_/X _1006_/Y _1013_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_39_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_641 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_836 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_858 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1136__C _1136_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_1_762 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1287__CLK _1294_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_36_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_749 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1486_ VGND VPWR _1486_/X _1486_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_933 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_977 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_counter.clk_A clkbuf_0_counter.clk/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1477 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0986__B _0993_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_110_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1805 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1271_ _1479_/A _1167_/Y _1271_/D _1279_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_96_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1351__264 la_data_out[42] _1351__264/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_209_333 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1789 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0986_ _1050_/B _0993_/D _0986_/Y _0999_/B _0986_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_140_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_693 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1302__CLK _1322_/CLK VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_173_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1057__B _1057_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_195_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1469_ VGND VPWR _1469_/X _1473_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_413 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1248__A _1248_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_137_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1335__248 io_out[35] _1335__248/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_144_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0840_ VGND VPWR _1503_/A _1505_/A _0840_/X _1502_/A _1504_/A VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_70_1241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0771_ VGND VPWR _0771_/X _0771_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0997__A _0997_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1323_ _1323_/Q _1258_/Y _1323_/D _1326_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_110_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1254_ VPWR VGND hold2/A _1254_/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1185_ VGND VPWR _1180_/X _1179_/X _1181_/X _1185_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_65_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1873 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0632__A1 _1503_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_833 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0969_ _0970_/B _0993_/D _0999_/B _0992_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_174_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput230 VPWR VGND wbs_dat_o[26] _0648_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_118_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1833 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput241 VPWR VGND wbs_dat_o[7] _0745_/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_160_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1877 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1421 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1793 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_794 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_777 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1561 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input62_A la_oenb[59] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_48_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1128__D _1142_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_174_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output149_A _1485_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_78_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1441__A _1473_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_130_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_917 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0823_ _0824_/A _0875_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1093 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_825 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0754_ VGND VPWR _1305_/D _0754_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_982 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_869 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0685_ VGND VPWR _1318_/D _0685_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1357__270 la_data_out[48] _1357__270/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_48_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1001 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1045 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1089 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1306_ _1306_/Q _1229_/Y _1306_/D _1322_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_97_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1785 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1237_ VGND VPWR _1231_/X _1230_/X _1232_/X _1237_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_84_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1168_ VPWR VGND _1203_/A hold2/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1099_ _1099_/A1 _0848_/X _1099_/Y _1143_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_53_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_731 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_797 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1925 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0908__A2 _0824_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_88_1365 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_357 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1393 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_637 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_569 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_961 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1449 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1861 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1171__A _1204_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1022_ _1022_/Y _0861_/X _1016_/B _0872_/B _1021_/X input77/X VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a311oi_4
XFILLER_130_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_497 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1821 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1805 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1849 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1589 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1049__C _1049_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_190_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0806_ _0838_/D _0922_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0737_ VGND VPWR _1308_/D _0737_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1901 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_0668_ VGND VPWR _0689_/S _1496_/A _1321_/Q _0669_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_118_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_861 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_937 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_609 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1645 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1017 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1373 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1009 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1033 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1077 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0934__A2_N _1497_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_120_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1061 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1256__A _1256_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_194_1777 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_97 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_922 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_955 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_454 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input25_A la_data_in[56] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_40_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_469 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_823 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_837 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_350 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1729 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1841 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1757 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1885 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1817 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1801 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_981 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1845 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1897 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1913 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1005_ VPWR VGND _1005_/X _1005_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_169_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1889 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1337 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_909 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1813 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1857 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1029 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_953 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1917 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0744__A0 _1481_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_103_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_881 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1869 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1073 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_553 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1057 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_973 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1505 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_697 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_809 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_949 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_853 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1085 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_993 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_897 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_525 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0983__B1 _0982_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_154_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_441 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1533 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_945 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_989 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_774 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_785 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1905 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_721 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1058__A4 _0832_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_781 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1649 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1037 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_829 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1673 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_841 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_385 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0974__B1 _0973_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_117_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_889 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1701 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1021 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1617 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1005 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1065 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1049 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1789 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_1485_ VGND VPWR _1485_/X _1485_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_797 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
.ends

